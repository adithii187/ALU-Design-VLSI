magic
tech scmos
magscale 9 1
timestamp 1700921468
<< nwell >>
rect 46 -126 67 -120
rect -6 -143 30 -133
rect 46 -138 63 -126
rect 46 -139 53 -138
rect 55 -139 63 -138
rect 46 -181 67 -175
rect -6 -198 30 -188
rect 46 -193 63 -181
rect 46 -194 53 -193
rect 55 -194 63 -193
rect 46 -227 67 -221
rect -6 -244 30 -234
rect 46 -239 63 -227
rect 46 -240 53 -239
rect 55 -240 63 -239
rect 46 -286 67 -280
rect -6 -303 30 -293
rect 46 -298 63 -286
rect 46 -299 53 -298
rect 55 -299 63 -298
rect 46 -339 67 -333
rect -6 -356 30 -346
rect 46 -351 63 -339
rect 46 -352 53 -351
rect 55 -352 63 -351
rect 46 -394 67 -388
rect -6 -411 30 -401
rect 46 -406 63 -394
rect 46 -407 53 -406
rect 55 -407 63 -406
rect 46 -440 67 -434
rect -6 -457 30 -447
rect 46 -452 63 -440
rect 46 -453 53 -452
rect 55 -453 63 -452
rect 46 -499 67 -493
rect -6 -516 30 -506
rect 46 -511 63 -499
rect 46 -512 53 -511
rect 55 -512 63 -511
<< ntransistor >>
rect 53 -148 55 -145
rect 2 -154 4 -151
rect 20 -154 22 -151
rect 53 -203 55 -200
rect 2 -209 4 -206
rect 20 -209 22 -206
rect 53 -249 55 -246
rect 2 -255 4 -252
rect 20 -255 22 -252
rect 53 -308 55 -305
rect 2 -314 4 -311
rect 20 -314 22 -311
rect 53 -361 55 -358
rect 2 -367 4 -364
rect 20 -367 22 -364
rect 53 -416 55 -413
rect 2 -422 4 -419
rect 20 -422 22 -419
rect 53 -462 55 -459
rect 2 -468 4 -465
rect 20 -468 22 -465
rect 53 -521 55 -518
rect 2 -527 4 -524
rect 20 -527 22 -524
<< ptransistor >>
rect 2 -140 4 -135
rect 20 -140 22 -135
rect 53 -137 55 -131
rect 2 -195 4 -190
rect 20 -195 22 -190
rect 53 -192 55 -186
rect 2 -241 4 -236
rect 20 -241 22 -236
rect 53 -238 55 -232
rect 2 -300 4 -295
rect 20 -300 22 -295
rect 53 -297 55 -291
rect 2 -353 4 -348
rect 20 -353 22 -348
rect 53 -350 55 -344
rect 2 -408 4 -403
rect 20 -408 22 -403
rect 53 -405 55 -399
rect 2 -454 4 -449
rect 20 -454 22 -449
rect 53 -451 55 -445
rect 2 -513 4 -508
rect 20 -513 22 -508
rect 53 -510 55 -504
<< ndiffusion >>
rect 48 -146 53 -145
rect 48 -148 49 -146
rect 52 -148 53 -146
rect 55 -148 57 -145
rect 60 -148 61 -145
rect -2 -152 2 -151
rect -2 -154 -1 -152
rect 1 -154 2 -152
rect 4 -154 20 -151
rect 22 -153 23 -151
rect 25 -153 26 -151
rect 22 -154 26 -153
rect 48 -201 53 -200
rect 48 -203 49 -201
rect 52 -203 53 -201
rect 55 -203 57 -200
rect 60 -203 61 -200
rect -2 -207 2 -206
rect -2 -209 -1 -207
rect 1 -209 2 -207
rect 4 -209 20 -206
rect 22 -208 23 -206
rect 25 -208 26 -206
rect 22 -209 26 -208
rect 48 -247 53 -246
rect 48 -249 49 -247
rect 52 -249 53 -247
rect 55 -249 57 -246
rect 60 -249 61 -246
rect -2 -253 2 -252
rect -2 -255 -1 -253
rect 1 -255 2 -253
rect 4 -255 20 -252
rect 22 -254 23 -252
rect 25 -254 26 -252
rect 22 -255 26 -254
rect 48 -306 53 -305
rect 48 -308 49 -306
rect 52 -308 53 -306
rect 55 -308 57 -305
rect 60 -308 61 -305
rect -2 -312 2 -311
rect -2 -314 -1 -312
rect 1 -314 2 -312
rect 4 -314 20 -311
rect 22 -313 23 -311
rect 25 -313 26 -311
rect 22 -314 26 -313
rect 48 -359 53 -358
rect 48 -361 49 -359
rect 52 -361 53 -359
rect 55 -361 57 -358
rect 60 -361 61 -358
rect -2 -365 2 -364
rect -2 -367 -1 -365
rect 1 -367 2 -365
rect 4 -367 20 -364
rect 22 -366 23 -364
rect 25 -366 26 -364
rect 22 -367 26 -366
rect 48 -414 53 -413
rect 48 -416 49 -414
rect 52 -416 53 -414
rect 55 -416 57 -413
rect 60 -416 61 -413
rect -2 -420 2 -419
rect -2 -422 -1 -420
rect 1 -422 2 -420
rect 4 -422 20 -419
rect 22 -421 23 -419
rect 25 -421 26 -419
rect 22 -422 26 -421
rect 48 -460 53 -459
rect 48 -462 49 -460
rect 52 -462 53 -460
rect 55 -462 57 -459
rect 60 -462 61 -459
rect -2 -466 2 -465
rect -2 -468 -1 -466
rect 1 -468 2 -466
rect 4 -468 20 -465
rect 22 -467 23 -465
rect 25 -467 26 -465
rect 22 -468 26 -467
rect 48 -519 53 -518
rect 48 -521 49 -519
rect 52 -521 53 -519
rect 55 -521 57 -518
rect 60 -521 61 -518
rect -2 -525 2 -524
rect -2 -527 -1 -525
rect 1 -527 2 -525
rect 4 -527 20 -524
rect 22 -526 23 -524
rect 25 -526 26 -524
rect 22 -527 26 -526
<< pdiffusion >>
rect 48 -134 49 -131
rect 52 -134 53 -131
rect -2 -136 2 -135
rect -2 -138 -1 -136
rect 1 -138 2 -136
rect -2 -140 2 -138
rect 4 -137 11 -135
rect 4 -139 5 -137
rect 7 -139 11 -137
rect 4 -140 11 -139
rect 15 -136 20 -135
rect 15 -138 16 -136
rect 18 -138 20 -136
rect 15 -140 20 -138
rect 22 -136 26 -135
rect 22 -138 23 -136
rect 25 -138 26 -136
rect 48 -137 53 -134
rect 55 -132 61 -131
rect 55 -135 57 -132
rect 60 -135 61 -132
rect 55 -137 61 -135
rect 22 -140 26 -138
rect 48 -189 49 -186
rect 52 -189 53 -186
rect -2 -191 2 -190
rect -2 -193 -1 -191
rect 1 -193 2 -191
rect -2 -195 2 -193
rect 4 -192 11 -190
rect 4 -194 5 -192
rect 7 -194 11 -192
rect 4 -195 11 -194
rect 15 -191 20 -190
rect 15 -193 16 -191
rect 18 -193 20 -191
rect 15 -195 20 -193
rect 22 -191 26 -190
rect 22 -193 23 -191
rect 25 -193 26 -191
rect 48 -192 53 -189
rect 55 -187 61 -186
rect 55 -190 57 -187
rect 60 -190 61 -187
rect 55 -192 61 -190
rect 22 -195 26 -193
rect 48 -235 49 -232
rect 52 -235 53 -232
rect -2 -237 2 -236
rect -2 -239 -1 -237
rect 1 -239 2 -237
rect -2 -241 2 -239
rect 4 -238 11 -236
rect 4 -240 5 -238
rect 7 -240 11 -238
rect 4 -241 11 -240
rect 15 -237 20 -236
rect 15 -239 16 -237
rect 18 -239 20 -237
rect 15 -241 20 -239
rect 22 -237 26 -236
rect 22 -239 23 -237
rect 25 -239 26 -237
rect 48 -238 53 -235
rect 55 -233 61 -232
rect 55 -236 57 -233
rect 60 -236 61 -233
rect 55 -238 61 -236
rect 22 -241 26 -239
rect 48 -294 49 -291
rect 52 -294 53 -291
rect -2 -296 2 -295
rect -2 -298 -1 -296
rect 1 -298 2 -296
rect -2 -300 2 -298
rect 4 -297 11 -295
rect 4 -299 5 -297
rect 7 -299 11 -297
rect 4 -300 11 -299
rect 15 -296 20 -295
rect 15 -298 16 -296
rect 18 -298 20 -296
rect 15 -300 20 -298
rect 22 -296 26 -295
rect 22 -298 23 -296
rect 25 -298 26 -296
rect 48 -297 53 -294
rect 55 -292 61 -291
rect 55 -295 57 -292
rect 60 -295 61 -292
rect 55 -297 61 -295
rect 22 -300 26 -298
rect 48 -347 49 -344
rect 52 -347 53 -344
rect -2 -349 2 -348
rect -2 -351 -1 -349
rect 1 -351 2 -349
rect -2 -353 2 -351
rect 4 -350 11 -348
rect 4 -352 5 -350
rect 7 -352 11 -350
rect 4 -353 11 -352
rect 15 -349 20 -348
rect 15 -351 16 -349
rect 18 -351 20 -349
rect 15 -353 20 -351
rect 22 -349 26 -348
rect 22 -351 23 -349
rect 25 -351 26 -349
rect 48 -350 53 -347
rect 55 -345 61 -344
rect 55 -348 57 -345
rect 60 -348 61 -345
rect 55 -350 61 -348
rect 22 -353 26 -351
rect 48 -402 49 -399
rect 52 -402 53 -399
rect -2 -404 2 -403
rect -2 -406 -1 -404
rect 1 -406 2 -404
rect -2 -408 2 -406
rect 4 -405 11 -403
rect 4 -407 5 -405
rect 7 -407 11 -405
rect 4 -408 11 -407
rect 15 -404 20 -403
rect 15 -406 16 -404
rect 18 -406 20 -404
rect 15 -408 20 -406
rect 22 -404 26 -403
rect 22 -406 23 -404
rect 25 -406 26 -404
rect 48 -405 53 -402
rect 55 -400 61 -399
rect 55 -403 57 -400
rect 60 -403 61 -400
rect 55 -405 61 -403
rect 22 -408 26 -406
rect 48 -448 49 -445
rect 52 -448 53 -445
rect -2 -450 2 -449
rect -2 -452 -1 -450
rect 1 -452 2 -450
rect -2 -454 2 -452
rect 4 -451 11 -449
rect 4 -453 5 -451
rect 7 -453 11 -451
rect 4 -454 11 -453
rect 15 -450 20 -449
rect 15 -452 16 -450
rect 18 -452 20 -450
rect 15 -454 20 -452
rect 22 -450 26 -449
rect 22 -452 23 -450
rect 25 -452 26 -450
rect 48 -451 53 -448
rect 55 -446 61 -445
rect 55 -449 57 -446
rect 60 -449 61 -446
rect 55 -451 61 -449
rect 22 -454 26 -452
rect 48 -507 49 -504
rect 52 -507 53 -504
rect -2 -509 2 -508
rect -2 -511 -1 -509
rect 1 -511 2 -509
rect -2 -513 2 -511
rect 4 -510 11 -508
rect 4 -512 5 -510
rect 7 -512 11 -510
rect 4 -513 11 -512
rect 15 -509 20 -508
rect 15 -511 16 -509
rect 18 -511 20 -509
rect 15 -513 20 -511
rect 22 -509 26 -508
rect 22 -511 23 -509
rect 25 -511 26 -509
rect 48 -510 53 -507
rect 55 -505 61 -504
rect 55 -508 57 -505
rect 60 -508 61 -505
rect 55 -510 61 -508
rect 22 -513 26 -511
<< ndcontact >>
rect 49 -149 52 -146
rect 57 -148 60 -145
rect -1 -154 1 -152
rect 23 -153 25 -151
rect 49 -204 52 -201
rect 57 -203 60 -200
rect -1 -209 1 -207
rect 23 -208 25 -206
rect 49 -250 52 -247
rect 57 -249 60 -246
rect -1 -255 1 -253
rect 23 -254 25 -252
rect 49 -309 52 -306
rect 57 -308 60 -305
rect -1 -314 1 -312
rect 23 -313 25 -311
rect 49 -362 52 -359
rect 57 -361 60 -358
rect -1 -367 1 -365
rect 23 -366 25 -364
rect 49 -417 52 -414
rect 57 -416 60 -413
rect -1 -422 1 -420
rect 23 -421 25 -419
rect 49 -463 52 -460
rect 57 -462 60 -459
rect -1 -468 1 -466
rect 23 -467 25 -465
rect 49 -522 52 -519
rect 57 -521 60 -518
rect -1 -527 1 -525
rect 23 -526 25 -524
<< pdcontact >>
rect 49 -134 52 -131
rect -1 -138 1 -136
rect 5 -139 7 -137
rect 16 -138 18 -136
rect 23 -138 25 -136
rect 57 -135 60 -132
rect 49 -189 52 -186
rect -1 -193 1 -191
rect 5 -194 7 -192
rect 16 -193 18 -191
rect 23 -193 25 -191
rect 57 -190 60 -187
rect 49 -235 52 -232
rect -1 -239 1 -237
rect 5 -240 7 -238
rect 16 -239 18 -237
rect 23 -239 25 -237
rect 57 -236 60 -233
rect 49 -294 52 -291
rect -1 -298 1 -296
rect 5 -299 7 -297
rect 16 -298 18 -296
rect 23 -298 25 -296
rect 57 -295 60 -292
rect 49 -347 52 -344
rect -1 -351 1 -349
rect 5 -352 7 -350
rect 16 -351 18 -349
rect 23 -351 25 -349
rect 57 -348 60 -345
rect 49 -402 52 -399
rect -1 -406 1 -404
rect 5 -407 7 -405
rect 16 -406 18 -404
rect 23 -406 25 -404
rect 57 -403 60 -400
rect 49 -448 52 -445
rect -1 -452 1 -450
rect 5 -453 7 -451
rect 16 -452 18 -450
rect 23 -452 25 -450
rect 57 -449 60 -446
rect 49 -507 52 -504
rect -1 -511 1 -509
rect 5 -512 7 -510
rect 16 -511 18 -509
rect 23 -511 25 -509
rect 57 -508 60 -505
<< polysilicon >>
rect 53 -131 55 -118
rect 2 -135 4 -132
rect 20 -135 22 -132
rect 2 -147 4 -140
rect -17 -149 4 -147
rect -17 -202 -15 -149
rect 2 -151 4 -149
rect 20 -151 22 -140
rect 53 -141 55 -137
rect 54 -144 55 -141
rect 53 -145 55 -144
rect 53 -150 55 -148
rect 2 -155 4 -154
rect 20 -155 22 -154
rect 53 -186 55 -173
rect 2 -190 4 -187
rect 20 -190 22 -187
rect 2 -202 4 -195
rect -17 -204 4 -202
rect -17 -249 -15 -204
rect 2 -206 4 -204
rect 20 -206 22 -195
rect 53 -196 55 -192
rect 54 -199 55 -196
rect 53 -200 55 -199
rect 53 -205 55 -203
rect 2 -210 4 -209
rect 20 -210 22 -209
rect 53 -232 55 -219
rect 2 -236 4 -233
rect 20 -236 22 -233
rect 2 -249 4 -241
rect -17 -251 4 -249
rect -17 -307 -15 -251
rect 2 -252 4 -251
rect 20 -252 22 -241
rect 53 -242 55 -238
rect 54 -245 55 -242
rect 53 -246 55 -245
rect 53 -251 55 -249
rect 2 -256 4 -255
rect 20 -256 22 -255
rect 53 -291 55 -278
rect 2 -295 4 -292
rect 20 -295 22 -292
rect 2 -307 4 -300
rect -17 -309 4 -307
rect -17 -360 -15 -309
rect 2 -311 4 -309
rect 20 -311 22 -300
rect 53 -301 55 -297
rect 54 -304 55 -301
rect 53 -305 55 -304
rect 53 -310 55 -308
rect 2 -315 4 -314
rect 20 -315 22 -314
rect 53 -344 55 -331
rect 2 -348 4 -345
rect 20 -348 22 -345
rect 2 -360 4 -353
rect -17 -362 4 -360
rect -17 -415 -15 -362
rect 2 -364 4 -362
rect 20 -364 22 -353
rect 53 -354 55 -350
rect 54 -357 55 -354
rect 53 -358 55 -357
rect 53 -363 55 -361
rect 2 -368 4 -367
rect 20 -368 22 -367
rect 53 -399 55 -386
rect 2 -403 4 -400
rect 20 -403 22 -400
rect 2 -415 4 -408
rect -17 -417 4 -415
rect -17 -462 -15 -417
rect 2 -419 4 -417
rect 20 -419 22 -408
rect 53 -409 55 -405
rect 54 -412 55 -409
rect 53 -413 55 -412
rect 53 -418 55 -416
rect 2 -423 4 -422
rect 20 -423 22 -422
rect 53 -445 55 -432
rect 2 -449 4 -446
rect 20 -449 22 -446
rect 2 -462 4 -454
rect -17 -464 4 -462
rect -17 -520 -15 -464
rect 2 -465 4 -464
rect 20 -465 22 -454
rect 53 -455 55 -451
rect 54 -458 55 -455
rect 53 -459 55 -458
rect 53 -464 55 -462
rect 2 -469 4 -468
rect 20 -469 22 -468
rect 53 -504 55 -491
rect 2 -508 4 -505
rect 20 -508 22 -505
rect 2 -520 4 -513
rect -17 -522 4 -520
rect 2 -524 4 -522
rect 20 -524 22 -513
rect 53 -514 55 -510
rect 54 -517 55 -514
rect 53 -518 55 -517
rect 53 -523 55 -521
rect 2 -528 4 -527
rect 20 -528 22 -527
<< polycontact >>
rect 51 -144 54 -141
rect 51 -199 54 -196
rect 51 -245 54 -242
rect 51 -304 54 -301
rect 51 -357 54 -354
rect 51 -412 54 -409
rect 51 -458 54 -455
rect 51 -517 54 -514
<< metal1 >>
rect 49 -125 76 -123
rect 49 -128 52 -125
rect -1 -130 52 -128
rect -1 -136 1 -130
rect 16 -136 18 -130
rect 49 -131 52 -130
rect 5 -145 7 -139
rect 23 -145 25 -138
rect 57 -140 60 -135
rect 41 -144 51 -141
rect 57 -143 63 -140
rect 41 -145 43 -144
rect 5 -147 43 -145
rect 57 -145 60 -143
rect 23 -151 25 -147
rect 49 -152 52 -149
rect -1 -156 1 -154
rect 49 -154 60 -152
rect 49 -156 53 -154
rect -13 -158 53 -156
rect -13 -211 -11 -158
rect 74 -178 76 -125
rect 49 -180 76 -178
rect 49 -183 52 -180
rect -1 -185 52 -183
rect -1 -191 1 -185
rect 16 -191 18 -185
rect 49 -186 52 -185
rect 5 -200 7 -194
rect 23 -200 25 -193
rect 57 -195 60 -190
rect 41 -199 51 -196
rect 57 -198 63 -195
rect 41 -200 43 -199
rect 5 -202 43 -200
rect 57 -200 60 -198
rect 23 -206 25 -202
rect 49 -207 52 -204
rect -1 -211 1 -209
rect 49 -209 60 -207
rect 49 -211 53 -209
rect -13 -213 53 -211
rect -13 -257 -11 -213
rect 74 -224 76 -180
rect 49 -226 76 -224
rect 49 -229 52 -226
rect -1 -231 52 -229
rect -1 -237 1 -231
rect 16 -237 18 -231
rect 49 -232 52 -231
rect 5 -246 7 -240
rect 23 -246 25 -239
rect 57 -241 60 -236
rect 41 -245 51 -242
rect 57 -244 63 -241
rect 41 -246 43 -245
rect 5 -248 43 -246
rect 57 -246 60 -244
rect 23 -252 25 -248
rect 49 -253 52 -250
rect -1 -257 1 -255
rect 49 -255 60 -253
rect 49 -257 53 -255
rect -13 -259 53 -257
rect -13 -316 -11 -259
rect 74 -283 76 -226
rect 49 -285 76 -283
rect 49 -288 52 -285
rect -1 -290 52 -288
rect -1 -296 1 -290
rect 16 -296 18 -290
rect 49 -291 52 -290
rect 5 -305 7 -299
rect 23 -305 25 -298
rect 57 -300 60 -295
rect 41 -304 51 -301
rect 57 -303 63 -300
rect 41 -305 43 -304
rect 5 -307 43 -305
rect 57 -305 60 -303
rect 23 -311 25 -307
rect 49 -312 52 -309
rect -1 -316 1 -314
rect 49 -314 60 -312
rect 49 -316 53 -314
rect -13 -318 53 -316
rect -13 -369 -11 -318
rect 74 -336 76 -285
rect 49 -338 76 -336
rect 49 -341 52 -338
rect -1 -343 52 -341
rect -1 -349 1 -343
rect 16 -349 18 -343
rect 49 -344 52 -343
rect 5 -358 7 -352
rect 23 -358 25 -351
rect 57 -353 60 -348
rect 41 -357 51 -354
rect 57 -356 63 -353
rect 41 -358 43 -357
rect 5 -360 43 -358
rect 57 -358 60 -356
rect 23 -364 25 -360
rect 49 -365 52 -362
rect -1 -369 1 -367
rect 49 -367 60 -365
rect 49 -369 53 -367
rect -13 -371 53 -369
rect -13 -424 -11 -371
rect 74 -391 76 -338
rect 49 -393 76 -391
rect 49 -396 52 -393
rect -1 -398 52 -396
rect -1 -404 1 -398
rect 16 -404 18 -398
rect 49 -399 52 -398
rect 5 -413 7 -407
rect 23 -413 25 -406
rect 57 -408 60 -403
rect 41 -412 51 -409
rect 57 -411 63 -408
rect 41 -413 43 -412
rect 5 -415 43 -413
rect 57 -413 60 -411
rect 23 -419 25 -415
rect 49 -420 52 -417
rect -1 -424 1 -422
rect 49 -422 60 -420
rect 49 -424 53 -422
rect -13 -426 53 -424
rect -13 -470 -11 -426
rect 74 -437 76 -393
rect 49 -439 76 -437
rect 49 -442 52 -439
rect -1 -444 52 -442
rect -1 -450 1 -444
rect 16 -450 18 -444
rect 49 -445 52 -444
rect 5 -459 7 -453
rect 23 -459 25 -452
rect 57 -454 60 -449
rect 41 -458 51 -455
rect 57 -457 63 -454
rect 41 -459 43 -458
rect 5 -461 43 -459
rect 57 -459 60 -457
rect 23 -465 25 -461
rect 49 -466 52 -463
rect -1 -470 1 -468
rect 49 -468 60 -466
rect 49 -470 53 -468
rect -13 -472 53 -470
rect -13 -529 -11 -472
rect 74 -496 76 -439
rect 49 -498 76 -496
rect 49 -501 52 -498
rect -1 -503 52 -501
rect -1 -509 1 -503
rect 16 -509 18 -503
rect 49 -504 52 -503
rect 5 -518 7 -512
rect 23 -518 25 -511
rect 57 -513 60 -508
rect 41 -517 51 -514
rect 57 -516 63 -513
rect 41 -518 43 -517
rect 5 -520 43 -518
rect 57 -518 60 -516
rect 23 -524 25 -520
rect 49 -525 52 -522
rect -1 -529 1 -527
rect 49 -527 60 -525
rect 49 -529 53 -527
rect -13 -531 53 -529
<< labels >>
rlabel polysilicon -16 -160 -16 -160 3 D2
rlabel polysilicon 21 -148 21 -148 1 a3
rlabel metal1 61 -142 61 -142 1 comp_a3
rlabel polysilicon 21 -204 21 -204 1 a2
rlabel metal1 61 -196 61 -196 1 comp_a2
rlabel polysilicon 21 -250 21 -250 1 a1
rlabel metal1 61 -242 61 -242 1 comp_a1
rlabel polysilicon 21 -309 21 -309 1 a0
rlabel metal1 61 -302 61 -302 1 comp_a0
rlabel polysilicon 21 -362 21 -362 1 b3
rlabel metal1 60 -355 60 -355 1 comp_b3
rlabel polysilicon 21 -416 21 -416 1 b2
rlabel metal1 61 -410 61 -410 1 comp_b2
rlabel polysilicon 21 -463 21 -463 1 b1
rlabel metal1 61 -455 61 -455 1 comp_b1
rlabel polysilicon 21 -522 21 -522 1 b0
rlabel metal1 61 -515 61 -515 1 comp_b0
rlabel metal1 75 -233 75 -233 7 vdd
rlabel metal1 -12 -239 -12 -239 3 gnd
<< end >>
