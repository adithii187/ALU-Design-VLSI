magic
tech scmos
timestamp 1700989981
<< nwell >>
rect 3141 4518 3249 5193
rect 3492 5121 3681 5166
rect 3501 5013 3654 5121
rect 3501 5004 3564 5013
rect 3582 5004 3654 5013
rect 3861 4815 4050 4860
rect 4707 4851 4896 4905
rect 3870 4707 4023 4815
rect 3870 4698 3933 4707
rect 3951 4698 4023 4707
rect 4239 4698 4563 4788
rect 4707 4743 4860 4851
rect 4707 4734 4770 4743
rect 4788 4734 4860 4743
rect 3141 3573 3249 4248
rect 3492 4176 3681 4221
rect 3501 4068 3654 4176
rect 3501 4059 3564 4068
rect 3582 4059 3654 4068
rect 3843 4023 4032 4050
rect 3834 4005 4032 4023
rect 4635 4041 4824 4095
rect 5463 4068 5652 4095
rect 5463 4050 5931 4068
rect 5463 4041 5652 4050
rect 3852 3897 4005 4005
rect 3852 3888 3915 3897
rect 3933 3888 4005 3897
rect 4167 3888 4491 3978
rect 4635 3933 4788 4041
rect 4635 3924 4698 3933
rect 4716 3924 4788 3933
rect 4995 3888 5319 3978
rect 5463 3933 5616 4041
rect 5913 4005 5931 4050
rect 5463 3924 5526 3933
rect 5544 3924 5616 3933
rect 5895 3888 6417 4005
rect 6201 3870 6237 3888
rect 4311 3249 5301 3276
rect 3141 2556 3249 3231
rect 4302 3222 5301 3249
rect 3492 3159 3672 3204
rect 3825 3159 4014 3204
rect 3501 3051 3654 3159
rect 3501 3042 3564 3051
rect 3582 3042 3654 3051
rect 3834 3051 3987 3159
rect 4311 3114 5301 3222
rect 3834 3042 3897 3051
rect 3915 3042 3987 3051
rect 4158 1953 5148 1980
rect 3141 1260 3249 1935
rect 4149 1926 5148 1953
rect 3492 1863 3672 1908
rect 3771 1863 3960 1908
rect 3501 1755 3654 1863
rect 3501 1746 3564 1755
rect 3582 1746 3654 1755
rect 3780 1755 3933 1863
rect 4158 1818 5148 1926
rect 3780 1746 3843 1755
rect 3861 1746 3933 1755
rect 3141 189 3249 864
rect 3492 792 3681 837
rect 3501 684 3654 792
rect 3501 675 3564 684
rect 3582 675 3654 684
rect 3861 486 4050 531
rect 4707 522 4896 576
rect 3870 378 4023 486
rect 3870 369 3933 378
rect 3951 369 4023 378
rect 4239 369 4563 459
rect 4707 414 4860 522
rect 4707 405 4770 414
rect 4788 405 4860 414
rect 3141 -756 3249 -81
rect 3492 -153 3681 -108
rect 3501 -261 3654 -153
rect 3501 -270 3564 -261
rect 3582 -270 3654 -261
rect 3843 -306 4032 -279
rect 3834 -324 4032 -306
rect 4635 -288 4824 -234
rect 5463 -261 5652 -234
rect 5463 -279 5931 -261
rect 5463 -288 5652 -279
rect 3852 -432 4005 -324
rect 3852 -441 3915 -432
rect 3933 -441 4005 -432
rect 4167 -441 4491 -351
rect 4635 -396 4788 -288
rect 4635 -405 4698 -396
rect 4716 -405 4788 -396
rect 4995 -441 5319 -351
rect 5463 -396 5616 -288
rect 5913 -324 5931 -279
rect 5463 -405 5526 -396
rect 5544 -405 5616 -396
rect 5895 -441 6417 -324
rect 6201 -459 6237 -441
rect 4311 -1080 5301 -1053
rect 3141 -1773 3249 -1098
rect 4302 -1107 5301 -1080
rect 3492 -1170 3672 -1125
rect 3825 -1170 4014 -1125
rect 3501 -1278 3654 -1170
rect 3501 -1287 3564 -1278
rect 3582 -1287 3654 -1278
rect 3834 -1278 3987 -1170
rect 4311 -1215 5301 -1107
rect 3834 -1287 3897 -1278
rect 3915 -1287 3987 -1278
rect 4158 -2376 5148 -2349
rect 3141 -3069 3249 -2394
rect 4149 -2403 5148 -2376
rect 3492 -2466 3672 -2421
rect 3771 -2466 3960 -2421
rect 3501 -2574 3654 -2466
rect 3501 -2583 3564 -2574
rect 3582 -2583 3654 -2574
rect 3780 -2574 3933 -2466
rect 4158 -2511 5148 -2403
rect 3780 -2583 3843 -2574
rect 3861 -2583 3933 -2574
rect 3141 -4608 3249 -3933
rect 3492 -4005 3681 -3960
rect 3501 -4113 3654 -4005
rect 3501 -4122 3564 -4113
rect 3582 -4122 3654 -4113
rect 3141 -5553 3249 -4878
rect 3492 -4950 3681 -4905
rect 3501 -5058 3654 -4950
rect 3501 -5067 3564 -5058
rect 3582 -5067 3654 -5058
rect 3141 -6570 3249 -5895
rect 3492 -5940 3681 -5922
rect 3699 -5940 3717 -4932
rect 4779 -5166 5769 -5004
rect 6606 -5013 6795 -4959
rect 6138 -5166 6462 -5076
rect 6606 -5121 6759 -5013
rect 6606 -5130 6669 -5121
rect 6687 -5130 6759 -5121
rect 3492 -5958 3717 -5940
rect 3492 -5967 3681 -5958
rect 3501 -6075 3654 -5967
rect 3501 -6084 3564 -6075
rect 3582 -6084 3654 -6075
rect 3141 -7866 3249 -7191
rect 3492 -7236 3681 -7218
rect 3699 -7236 3717 -5958
rect 3492 -7254 3717 -7236
rect 3492 -7263 3681 -7254
rect 3501 -7371 3654 -7263
rect 3501 -7380 3564 -7371
rect 3582 -7380 3654 -7371
<< ntransistor >>
rect 2916 5112 2970 5130
rect 2916 4941 2970 4959
rect 3564 4923 3582 4950
rect 2916 4743 2970 4761
rect 2916 4581 2970 4599
rect 3933 4617 3951 4644
rect 4770 4653 4788 4680
rect 4311 4599 4329 4626
rect 4419 4599 4428 4626
rect 4473 4599 4491 4626
rect 2916 4167 2970 4185
rect 2916 3996 2970 4014
rect 3564 3978 3582 4005
rect 2916 3798 2970 3816
rect 3915 3807 3933 3834
rect 4698 3843 4716 3870
rect 5526 3843 5544 3870
rect 4239 3789 4257 3816
rect 4347 3789 4356 3816
rect 4401 3789 4419 3816
rect 5067 3789 5085 3816
rect 5229 3789 5247 3816
rect 5949 3789 5967 3816
rect 6039 3789 6057 3816
rect 6129 3789 6147 3816
rect 6219 3789 6237 3816
rect 6345 3789 6363 3816
rect 2916 3636 2970 3654
rect 2916 3150 2970 3168
rect 2916 2979 2970 2997
rect 3564 2961 3582 2988
rect 3897 2961 3915 2988
rect 4401 2979 4419 3006
rect 4527 2979 4545 3006
rect 4671 2979 4689 3006
rect 4797 2979 4815 3006
rect 4932 2979 4950 3006
rect 5193 2979 5211 3006
rect 2916 2781 2970 2799
rect 2916 2619 2970 2637
rect 2916 1854 2970 1872
rect 2916 1683 2970 1701
rect 3564 1665 3582 1692
rect 3843 1665 3861 1692
rect 4248 1683 4266 1710
rect 4374 1683 4392 1710
rect 4518 1683 4536 1710
rect 4644 1683 4662 1710
rect 4779 1683 4797 1710
rect 5040 1683 5058 1710
rect 2916 1485 2970 1503
rect 2916 1323 2970 1341
rect 2916 783 2970 801
rect 2916 612 2970 630
rect 3564 594 3582 621
rect 2916 414 2970 432
rect 2916 252 2970 270
rect 3933 288 3951 315
rect 4770 324 4788 351
rect 4311 270 4329 297
rect 4419 270 4428 297
rect 4473 270 4491 297
rect 2916 -162 2970 -144
rect 2916 -333 2970 -315
rect 3564 -351 3582 -324
rect 2916 -531 2970 -513
rect 3915 -522 3933 -495
rect 4698 -486 4716 -459
rect 5526 -486 5544 -459
rect 4239 -540 4257 -513
rect 4347 -540 4356 -513
rect 4401 -540 4419 -513
rect 5067 -540 5085 -513
rect 5229 -540 5247 -513
rect 5949 -540 5967 -513
rect 6039 -540 6057 -513
rect 6129 -540 6147 -513
rect 6219 -540 6237 -513
rect 6345 -540 6363 -513
rect 2916 -693 2970 -675
rect 2916 -1179 2970 -1161
rect 2916 -1350 2970 -1332
rect 3564 -1368 3582 -1341
rect 3897 -1368 3915 -1341
rect 4401 -1350 4419 -1323
rect 4527 -1350 4545 -1323
rect 4671 -1350 4689 -1323
rect 4797 -1350 4815 -1323
rect 4932 -1350 4950 -1323
rect 5193 -1350 5211 -1323
rect 2916 -1548 2970 -1530
rect 2916 -1710 2970 -1692
rect 2916 -2475 2970 -2457
rect 2916 -2646 2970 -2628
rect 3564 -2664 3582 -2637
rect 2916 -2844 2970 -2826
rect 2916 -3006 2970 -2988
rect 2916 -4014 2970 -3996
rect 3843 -2664 3861 -2637
rect 4248 -2646 4266 -2619
rect 4374 -2646 4392 -2619
rect 4518 -2646 4536 -2619
rect 4644 -2646 4662 -2619
rect 4779 -2646 4797 -2619
rect 5040 -2646 5058 -2619
rect 2916 -4185 2970 -4167
rect 3564 -4203 3582 -4176
rect 2916 -4383 2970 -4365
rect 2916 -4545 2970 -4527
rect 2916 -4959 2970 -4941
rect 2916 -5130 2970 -5112
rect 3564 -5148 3582 -5121
rect 2916 -5328 2970 -5310
rect 6669 -5211 6687 -5184
rect 6210 -5265 6228 -5238
rect 6372 -5265 6390 -5238
rect 4869 -5301 4887 -5274
rect 4995 -5301 5013 -5274
rect 5139 -5301 5157 -5274
rect 5265 -5301 5283 -5274
rect 5400 -5301 5418 -5274
rect 5661 -5301 5679 -5274
rect 2916 -5490 2970 -5472
rect 2916 -5976 2970 -5958
rect 2916 -6147 2970 -6129
rect 3564 -6165 3582 -6138
rect 2916 -6345 2970 -6327
rect 2916 -6507 2970 -6489
rect 2916 -7272 2970 -7254
rect 2916 -7443 2970 -7425
rect 3564 -7461 3582 -7434
rect 2916 -7641 2970 -7623
rect 2916 -7803 2970 -7785
<< ptransistor >>
rect 3168 5112 3231 5130
rect 3564 5022 3582 5076
rect 3168 4941 3231 4959
rect 3168 4743 3231 4761
rect 3168 4581 3231 4599
rect 3933 4716 3951 4770
rect 4311 4725 4329 4770
rect 4473 4725 4491 4770
rect 4770 4752 4788 4806
rect 3168 4167 3231 4185
rect 3564 4077 3582 4131
rect 3168 3996 3231 4014
rect 3168 3798 3231 3816
rect 3915 3906 3933 3960
rect 4239 3915 4257 3960
rect 4401 3915 4419 3960
rect 4698 3942 4716 3996
rect 5067 3915 5085 3960
rect 5229 3915 5247 3960
rect 5526 3942 5544 3996
rect 5949 3906 5967 3951
rect 6003 3906 6021 3951
rect 6039 3906 6057 3951
rect 6129 3906 6147 3951
rect 6219 3906 6237 3951
rect 6345 3906 6363 3951
rect 3168 3636 3231 3654
rect 3168 3150 3231 3168
rect 4401 3132 4419 3186
rect 4527 3132 4545 3186
rect 4671 3132 4689 3186
rect 4797 3132 4815 3186
rect 4932 3132 4950 3186
rect 5193 3132 5211 3186
rect 3564 3060 3582 3114
rect 3897 3060 3915 3114
rect 3168 2979 3231 2997
rect 3168 2781 3231 2799
rect 3168 2619 3231 2637
rect 3168 1854 3231 1872
rect 4248 1836 4266 1890
rect 4374 1836 4392 1890
rect 4518 1836 4536 1890
rect 4644 1836 4662 1890
rect 4779 1836 4797 1890
rect 5040 1836 5058 1890
rect 3564 1764 3582 1818
rect 3843 1764 3861 1818
rect 3168 1683 3231 1701
rect 3168 1485 3231 1503
rect 3168 1323 3231 1341
rect 3168 783 3231 801
rect 3564 693 3582 747
rect 3168 612 3231 630
rect 3168 414 3231 432
rect 3168 252 3231 270
rect 3933 387 3951 441
rect 4311 396 4329 441
rect 4473 396 4491 441
rect 4770 423 4788 477
rect 3168 -162 3231 -144
rect 3564 -252 3582 -198
rect 3168 -333 3231 -315
rect 3168 -531 3231 -513
rect 3915 -423 3933 -369
rect 4239 -414 4257 -369
rect 4401 -414 4419 -369
rect 4698 -387 4716 -333
rect 5067 -414 5085 -369
rect 5229 -414 5247 -369
rect 5526 -387 5544 -333
rect 5949 -423 5967 -378
rect 6003 -423 6021 -378
rect 6039 -423 6057 -378
rect 6129 -423 6147 -378
rect 6219 -423 6237 -378
rect 6345 -423 6363 -378
rect 3168 -693 3231 -675
rect 3168 -1179 3231 -1161
rect 4401 -1197 4419 -1143
rect 4527 -1197 4545 -1143
rect 4671 -1197 4689 -1143
rect 4797 -1197 4815 -1143
rect 4932 -1197 4950 -1143
rect 5193 -1197 5211 -1143
rect 3564 -1269 3582 -1215
rect 3897 -1269 3915 -1215
rect 3168 -1350 3231 -1332
rect 3168 -1548 3231 -1530
rect 3168 -1710 3231 -1692
rect 3168 -2475 3231 -2457
rect 3564 -2565 3582 -2511
rect 3168 -2646 3231 -2628
rect 3168 -2844 3231 -2826
rect 3168 -3006 3231 -2988
rect 3168 -4014 3231 -3996
rect 4248 -2493 4266 -2439
rect 4374 -2493 4392 -2439
rect 4518 -2493 4536 -2439
rect 4644 -2493 4662 -2439
rect 4779 -2493 4797 -2439
rect 5040 -2493 5058 -2439
rect 3843 -2565 3861 -2511
rect 3564 -4104 3582 -4050
rect 3168 -4185 3231 -4167
rect 3168 -4383 3231 -4365
rect 3168 -4545 3231 -4527
rect 3168 -4959 3231 -4941
rect 3564 -5049 3582 -4995
rect 3168 -5130 3231 -5112
rect 3168 -5328 3231 -5310
rect 4869 -5148 4887 -5094
rect 4995 -5148 5013 -5094
rect 5139 -5148 5157 -5094
rect 5265 -5148 5283 -5094
rect 5400 -5148 5418 -5094
rect 5661 -5148 5679 -5094
rect 6210 -5139 6228 -5094
rect 6372 -5139 6390 -5094
rect 6669 -5112 6687 -5058
rect 3168 -5490 3231 -5472
rect 3168 -5976 3231 -5958
rect 3564 -6066 3582 -6012
rect 3168 -6147 3231 -6129
rect 3168 -6345 3231 -6327
rect 3168 -6507 3231 -6489
rect 3168 -7272 3231 -7254
rect 3564 -7362 3582 -7308
rect 3168 -7443 3231 -7425
rect 3168 -7641 3231 -7623
rect 3168 -7803 3231 -7785
<< ndiffusion >>
rect 2916 5175 2970 5184
rect 2916 5139 2925 5175
rect 2961 5139 2970 5175
rect 2916 5130 2970 5139
rect 2916 5103 2970 5112
rect 2916 5067 2925 5103
rect 2961 5067 2970 5103
rect 2916 5058 2970 5067
rect 2916 5004 2970 5013
rect 2916 4968 2925 5004
rect 2961 4968 2970 5004
rect 2916 4959 2970 4968
rect 3519 4941 3564 4950
rect 2916 4932 2970 4941
rect 2916 4896 2925 4932
rect 2961 4896 2970 4932
rect 2916 4887 2970 4896
rect 3519 4923 3528 4941
rect 3555 4923 3564 4941
rect 3582 4923 3600 4950
rect 3627 4923 3636 4950
rect 2916 4815 2970 4824
rect 2916 4779 2925 4815
rect 2961 4779 2970 4815
rect 2916 4761 2970 4779
rect 2916 4734 2970 4743
rect 2916 4698 2925 4734
rect 2961 4698 2970 4734
rect 2916 4689 2970 4698
rect 2916 4653 2970 4662
rect 2916 4617 2925 4653
rect 2961 4617 2970 4653
rect 2916 4599 2970 4617
rect 2916 4572 2970 4581
rect 2916 4536 2925 4572
rect 2961 4536 2970 4572
rect 2916 4527 2970 4536
rect 3888 4635 3933 4644
rect 3888 4617 3897 4635
rect 3924 4617 3933 4635
rect 3951 4617 3969 4644
rect 3996 4617 4005 4644
rect 4725 4671 4770 4680
rect 4725 4653 4734 4671
rect 4761 4653 4770 4671
rect 4788 4653 4806 4680
rect 4833 4653 4842 4680
rect 4275 4617 4311 4626
rect 4275 4599 4284 4617
rect 4302 4599 4311 4617
rect 4329 4599 4419 4626
rect 4428 4599 4473 4626
rect 4491 4608 4500 4626
rect 4518 4608 4527 4626
rect 4491 4599 4527 4608
rect 2916 4230 2970 4239
rect 2916 4194 2925 4230
rect 2961 4194 2970 4230
rect 2916 4185 2970 4194
rect 2916 4158 2970 4167
rect 2916 4122 2925 4158
rect 2961 4122 2970 4158
rect 2916 4113 2970 4122
rect 2916 4059 2970 4068
rect 2916 4023 2925 4059
rect 2961 4023 2970 4059
rect 2916 4014 2970 4023
rect 3519 3996 3564 4005
rect 2916 3987 2970 3996
rect 2916 3951 2925 3987
rect 2961 3951 2970 3987
rect 2916 3942 2970 3951
rect 3519 3978 3528 3996
rect 3555 3978 3564 3996
rect 3582 3978 3600 4005
rect 3627 3978 3636 4005
rect 2916 3870 2970 3879
rect 2916 3834 2925 3870
rect 2961 3834 2970 3870
rect 2916 3816 2970 3834
rect 2916 3789 2970 3798
rect 2916 3753 2925 3789
rect 2961 3753 2970 3789
rect 2916 3744 2970 3753
rect 3870 3825 3915 3834
rect 3870 3807 3879 3825
rect 3906 3807 3915 3825
rect 3933 3807 3951 3834
rect 3978 3807 3987 3834
rect 4653 3861 4698 3870
rect 4653 3843 4662 3861
rect 4689 3843 4698 3861
rect 4716 3843 4734 3870
rect 4761 3843 4770 3870
rect 5481 3861 5526 3870
rect 5481 3843 5490 3861
rect 5517 3843 5526 3861
rect 5544 3843 5562 3870
rect 5589 3843 5598 3870
rect 4203 3807 4239 3816
rect 4203 3789 4212 3807
rect 4230 3789 4239 3807
rect 4257 3789 4347 3816
rect 4356 3789 4401 3816
rect 4419 3798 4428 3816
rect 4446 3798 4455 3816
rect 4419 3789 4455 3798
rect 5031 3807 5067 3816
rect 5031 3789 5040 3807
rect 5058 3789 5067 3807
rect 5085 3789 5229 3816
rect 5247 3798 5256 3816
rect 5274 3798 5283 3816
rect 5247 3789 5283 3798
rect 5904 3798 5913 3816
rect 5931 3798 5949 3816
rect 5904 3789 5949 3798
rect 5967 3798 5976 3816
rect 5967 3789 5994 3798
rect 6003 3798 6012 3816
rect 6030 3798 6039 3816
rect 6003 3789 6039 3798
rect 6057 3798 6066 3816
rect 6057 3789 6084 3798
rect 6093 3798 6102 3816
rect 6120 3798 6129 3816
rect 6093 3789 6129 3798
rect 6147 3798 6156 3816
rect 6147 3789 6174 3798
rect 6183 3798 6192 3816
rect 6210 3798 6219 3816
rect 6183 3789 6219 3798
rect 6237 3798 6246 3816
rect 6237 3789 6264 3798
rect 6309 3798 6318 3816
rect 6336 3798 6345 3816
rect 6309 3789 6345 3798
rect 6363 3798 6372 3816
rect 6390 3798 6399 3816
rect 6363 3789 6399 3798
rect 2916 3708 2970 3717
rect 2916 3672 2925 3708
rect 2961 3672 2970 3708
rect 2916 3654 2970 3672
rect 2916 3627 2970 3636
rect 2916 3591 2925 3627
rect 2961 3591 2970 3627
rect 2916 3582 2970 3591
rect 2916 3213 2970 3222
rect 2916 3177 2925 3213
rect 2961 3177 2970 3213
rect 2916 3168 2970 3177
rect 2916 3141 2970 3150
rect 2916 3105 2925 3141
rect 2961 3105 2970 3141
rect 2916 3096 2970 3105
rect 2916 3042 2970 3051
rect 2916 3006 2925 3042
rect 2961 3006 2970 3042
rect 2916 2997 2970 3006
rect 3519 2979 3564 2988
rect 2916 2970 2970 2979
rect 2916 2934 2925 2970
rect 2961 2934 2970 2970
rect 2916 2925 2970 2934
rect 3519 2961 3528 2979
rect 3555 2961 3564 2979
rect 3582 2961 3600 2988
rect 3627 2961 3636 2988
rect 3852 2979 3897 2988
rect 3852 2961 3861 2979
rect 3888 2961 3897 2979
rect 3915 2961 3933 2988
rect 3960 2961 3969 2988
rect 4356 2979 4365 3006
rect 4392 2979 4401 3006
rect 4419 2979 4527 3006
rect 4545 2979 4671 3006
rect 4689 2979 4797 3006
rect 4815 2979 4932 3006
rect 4950 2979 4986 3006
rect 5013 2979 5085 3006
rect 5139 2979 5157 3006
rect 5184 2979 5193 3006
rect 5211 2979 5220 3006
rect 5247 2979 5256 3006
rect 2916 2853 2970 2862
rect 2916 2817 2925 2853
rect 2961 2817 2970 2853
rect 2916 2799 2970 2817
rect 2916 2772 2970 2781
rect 2916 2736 2925 2772
rect 2961 2736 2970 2772
rect 2916 2727 2970 2736
rect 2916 2691 2970 2700
rect 2916 2655 2925 2691
rect 2961 2655 2970 2691
rect 2916 2637 2970 2655
rect 2916 2610 2970 2619
rect 2916 2574 2925 2610
rect 2961 2574 2970 2610
rect 2916 2565 2970 2574
rect 2916 1917 2970 1926
rect 2916 1881 2925 1917
rect 2961 1881 2970 1917
rect 2916 1872 2970 1881
rect 2916 1845 2970 1854
rect 2916 1809 2925 1845
rect 2961 1809 2970 1845
rect 2916 1800 2970 1809
rect 2916 1746 2970 1755
rect 2916 1710 2925 1746
rect 2961 1710 2970 1746
rect 2916 1701 2970 1710
rect 3519 1683 3564 1692
rect 2916 1674 2970 1683
rect 2916 1638 2925 1674
rect 2961 1638 2970 1674
rect 2916 1629 2970 1638
rect 3519 1665 3528 1683
rect 3555 1665 3564 1683
rect 3582 1665 3600 1692
rect 3627 1665 3636 1692
rect 3798 1683 3843 1692
rect 3798 1665 3807 1683
rect 3834 1665 3843 1683
rect 3861 1665 3879 1692
rect 3906 1665 3915 1692
rect 4203 1683 4212 1710
rect 4239 1683 4248 1710
rect 4266 1683 4374 1710
rect 4392 1683 4518 1710
rect 4536 1683 4644 1710
rect 4662 1683 4779 1710
rect 4797 1683 4833 1710
rect 4860 1683 4932 1710
rect 4986 1683 5004 1710
rect 5031 1683 5040 1710
rect 5058 1683 5067 1710
rect 5094 1683 5103 1710
rect 2916 1557 2970 1566
rect 2916 1521 2925 1557
rect 2961 1521 2970 1557
rect 2916 1503 2970 1521
rect 2916 1476 2970 1485
rect 2916 1440 2925 1476
rect 2961 1440 2970 1476
rect 2916 1431 2970 1440
rect 2916 1395 2970 1404
rect 2916 1359 2925 1395
rect 2961 1359 2970 1395
rect 2916 1341 2970 1359
rect 2916 1314 2970 1323
rect 2916 1278 2925 1314
rect 2961 1278 2970 1314
rect 2916 1269 2970 1278
rect 2916 846 2970 855
rect 2916 810 2925 846
rect 2961 810 2970 846
rect 2916 801 2970 810
rect 2916 774 2970 783
rect 2916 738 2925 774
rect 2961 738 2970 774
rect 2916 729 2970 738
rect 2916 675 2970 684
rect 2916 639 2925 675
rect 2961 639 2970 675
rect 2916 630 2970 639
rect 3519 612 3564 621
rect 2916 603 2970 612
rect 2916 567 2925 603
rect 2961 567 2970 603
rect 2916 558 2970 567
rect 3519 594 3528 612
rect 3555 594 3564 612
rect 3582 594 3600 621
rect 3627 594 3636 621
rect 2916 486 2970 495
rect 2916 450 2925 486
rect 2961 450 2970 486
rect 2916 432 2970 450
rect 2916 405 2970 414
rect 2916 369 2925 405
rect 2961 369 2970 405
rect 2916 360 2970 369
rect 2916 324 2970 333
rect 2916 288 2925 324
rect 2961 288 2970 324
rect 2916 270 2970 288
rect 2916 243 2970 252
rect 2916 207 2925 243
rect 2961 207 2970 243
rect 2916 198 2970 207
rect 3888 306 3933 315
rect 3888 288 3897 306
rect 3924 288 3933 306
rect 3951 288 3969 315
rect 3996 288 4005 315
rect 4725 342 4770 351
rect 4725 324 4734 342
rect 4761 324 4770 342
rect 4788 324 4806 351
rect 4833 324 4842 351
rect 4275 288 4311 297
rect 4275 270 4284 288
rect 4302 270 4311 288
rect 4329 270 4419 297
rect 4428 270 4473 297
rect 4491 279 4500 297
rect 4518 279 4527 297
rect 4491 270 4527 279
rect 2916 -99 2970 -90
rect 2916 -135 2925 -99
rect 2961 -135 2970 -99
rect 2916 -144 2970 -135
rect 2916 -171 2970 -162
rect 2916 -207 2925 -171
rect 2961 -207 2970 -171
rect 2916 -216 2970 -207
rect 2916 -270 2970 -261
rect 2916 -306 2925 -270
rect 2961 -306 2970 -270
rect 2916 -315 2970 -306
rect 3519 -333 3564 -324
rect 2916 -342 2970 -333
rect 2916 -378 2925 -342
rect 2961 -378 2970 -342
rect 2916 -387 2970 -378
rect 3519 -351 3528 -333
rect 3555 -351 3564 -333
rect 3582 -351 3600 -324
rect 3627 -351 3636 -324
rect 2916 -459 2970 -450
rect 2916 -495 2925 -459
rect 2961 -495 2970 -459
rect 2916 -513 2970 -495
rect 2916 -540 2970 -531
rect 2916 -576 2925 -540
rect 2961 -576 2970 -540
rect 2916 -585 2970 -576
rect 3870 -504 3915 -495
rect 3870 -522 3879 -504
rect 3906 -522 3915 -504
rect 3933 -522 3951 -495
rect 3978 -522 3987 -495
rect 4653 -468 4698 -459
rect 4653 -486 4662 -468
rect 4689 -486 4698 -468
rect 4716 -486 4734 -459
rect 4761 -486 4770 -459
rect 5481 -468 5526 -459
rect 5481 -486 5490 -468
rect 5517 -486 5526 -468
rect 5544 -486 5562 -459
rect 5589 -486 5598 -459
rect 4203 -522 4239 -513
rect 4203 -540 4212 -522
rect 4230 -540 4239 -522
rect 4257 -540 4347 -513
rect 4356 -540 4401 -513
rect 4419 -531 4428 -513
rect 4446 -531 4455 -513
rect 4419 -540 4455 -531
rect 5031 -522 5067 -513
rect 5031 -540 5040 -522
rect 5058 -540 5067 -522
rect 5085 -540 5229 -513
rect 5247 -531 5256 -513
rect 5274 -531 5283 -513
rect 5247 -540 5283 -531
rect 5904 -531 5913 -513
rect 5931 -531 5949 -513
rect 5904 -540 5949 -531
rect 5967 -531 5976 -513
rect 5967 -540 5994 -531
rect 6003 -531 6012 -513
rect 6030 -531 6039 -513
rect 6003 -540 6039 -531
rect 6057 -531 6066 -513
rect 6057 -540 6084 -531
rect 6093 -531 6102 -513
rect 6120 -531 6129 -513
rect 6093 -540 6129 -531
rect 6147 -531 6156 -513
rect 6147 -540 6174 -531
rect 6183 -531 6192 -513
rect 6210 -531 6219 -513
rect 6183 -540 6219 -531
rect 6237 -531 6246 -513
rect 6237 -540 6264 -531
rect 6309 -531 6318 -513
rect 6336 -531 6345 -513
rect 6309 -540 6345 -531
rect 6363 -531 6372 -513
rect 6390 -531 6399 -513
rect 6363 -540 6399 -531
rect 2916 -621 2970 -612
rect 2916 -657 2925 -621
rect 2961 -657 2970 -621
rect 2916 -675 2970 -657
rect 2916 -702 2970 -693
rect 2916 -738 2925 -702
rect 2961 -738 2970 -702
rect 2916 -747 2970 -738
rect 2916 -1116 2970 -1107
rect 2916 -1152 2925 -1116
rect 2961 -1152 2970 -1116
rect 2916 -1161 2970 -1152
rect 2916 -1188 2970 -1179
rect 2916 -1224 2925 -1188
rect 2961 -1224 2970 -1188
rect 2916 -1233 2970 -1224
rect 2916 -1287 2970 -1278
rect 2916 -1323 2925 -1287
rect 2961 -1323 2970 -1287
rect 2916 -1332 2970 -1323
rect 3519 -1350 3564 -1341
rect 2916 -1359 2970 -1350
rect 2916 -1395 2925 -1359
rect 2961 -1395 2970 -1359
rect 2916 -1404 2970 -1395
rect 3519 -1368 3528 -1350
rect 3555 -1368 3564 -1350
rect 3582 -1368 3600 -1341
rect 3627 -1368 3636 -1341
rect 3852 -1350 3897 -1341
rect 3852 -1368 3861 -1350
rect 3888 -1368 3897 -1350
rect 3915 -1368 3933 -1341
rect 3960 -1368 3969 -1341
rect 4356 -1350 4365 -1323
rect 4392 -1350 4401 -1323
rect 4419 -1350 4527 -1323
rect 4545 -1350 4671 -1323
rect 4689 -1350 4797 -1323
rect 4815 -1350 4932 -1323
rect 4950 -1350 4986 -1323
rect 5013 -1350 5085 -1323
rect 5139 -1350 5157 -1323
rect 5184 -1350 5193 -1323
rect 5211 -1350 5220 -1323
rect 5247 -1350 5256 -1323
rect 2916 -1476 2970 -1467
rect 2916 -1512 2925 -1476
rect 2961 -1512 2970 -1476
rect 2916 -1530 2970 -1512
rect 2916 -1557 2970 -1548
rect 2916 -1593 2925 -1557
rect 2961 -1593 2970 -1557
rect 2916 -1602 2970 -1593
rect 2916 -1638 2970 -1629
rect 2916 -1674 2925 -1638
rect 2961 -1674 2970 -1638
rect 2916 -1692 2970 -1674
rect 2916 -1719 2970 -1710
rect 2916 -1755 2925 -1719
rect 2961 -1755 2970 -1719
rect 2916 -1764 2970 -1755
rect 2916 -2412 2970 -2403
rect 2916 -2448 2925 -2412
rect 2961 -2448 2970 -2412
rect 2916 -2457 2970 -2448
rect 2916 -2484 2970 -2475
rect 2916 -2520 2925 -2484
rect 2961 -2520 2970 -2484
rect 2916 -2529 2970 -2520
rect 2916 -2583 2970 -2574
rect 2916 -2619 2925 -2583
rect 2961 -2619 2970 -2583
rect 2916 -2628 2970 -2619
rect 3519 -2646 3564 -2637
rect 2916 -2655 2970 -2646
rect 2916 -2691 2925 -2655
rect 2961 -2691 2970 -2655
rect 2916 -2700 2970 -2691
rect 3519 -2664 3528 -2646
rect 3555 -2664 3564 -2646
rect 3582 -2664 3600 -2637
rect 3627 -2664 3636 -2637
rect 2916 -2772 2970 -2763
rect 2916 -2808 2925 -2772
rect 2961 -2808 2970 -2772
rect 2916 -2826 2970 -2808
rect 2916 -2853 2970 -2844
rect 2916 -2889 2925 -2853
rect 2961 -2889 2970 -2853
rect 2916 -2898 2970 -2889
rect 2916 -2934 2970 -2925
rect 2916 -2970 2925 -2934
rect 2961 -2970 2970 -2934
rect 2916 -2988 2970 -2970
rect 2916 -3015 2970 -3006
rect 2916 -3051 2925 -3015
rect 2961 -3051 2970 -3015
rect 2916 -3060 2970 -3051
rect 2916 -3951 2970 -3942
rect 2916 -3987 2925 -3951
rect 2961 -3987 2970 -3951
rect 2916 -3996 2970 -3987
rect 2916 -4023 2970 -4014
rect 2916 -4059 2925 -4023
rect 2961 -4059 2970 -4023
rect 2916 -4068 2970 -4059
rect 2916 -4122 2970 -4113
rect 2916 -4158 2925 -4122
rect 2961 -4158 2970 -4122
rect 2916 -4167 2970 -4158
rect 3798 -2646 3843 -2637
rect 3798 -2664 3807 -2646
rect 3834 -2664 3843 -2646
rect 3861 -2664 3879 -2637
rect 3906 -2664 3915 -2637
rect 4203 -2646 4212 -2619
rect 4239 -2646 4248 -2619
rect 4266 -2646 4374 -2619
rect 4392 -2646 4518 -2619
rect 4536 -2646 4644 -2619
rect 4662 -2646 4779 -2619
rect 4797 -2646 4833 -2619
rect 4860 -2646 4932 -2619
rect 4986 -2646 5004 -2619
rect 5031 -2646 5040 -2619
rect 5058 -2646 5067 -2619
rect 5094 -2646 5103 -2619
rect 3519 -4185 3564 -4176
rect 2916 -4194 2970 -4185
rect 2916 -4230 2925 -4194
rect 2961 -4230 2970 -4194
rect 2916 -4239 2970 -4230
rect 3519 -4203 3528 -4185
rect 3555 -4203 3564 -4185
rect 3582 -4203 3600 -4176
rect 3627 -4203 3636 -4176
rect 2916 -4311 2970 -4302
rect 2916 -4347 2925 -4311
rect 2961 -4347 2970 -4311
rect 2916 -4365 2970 -4347
rect 2916 -4392 2970 -4383
rect 2916 -4428 2925 -4392
rect 2961 -4428 2970 -4392
rect 2916 -4437 2970 -4428
rect 2916 -4473 2970 -4464
rect 2916 -4509 2925 -4473
rect 2961 -4509 2970 -4473
rect 2916 -4527 2970 -4509
rect 2916 -4554 2970 -4545
rect 2916 -4590 2925 -4554
rect 2961 -4590 2970 -4554
rect 2916 -4599 2970 -4590
rect 2916 -4896 2970 -4887
rect 2916 -4932 2925 -4896
rect 2961 -4932 2970 -4896
rect 2916 -4941 2970 -4932
rect 2916 -4968 2970 -4959
rect 2916 -5004 2925 -4968
rect 2961 -5004 2970 -4968
rect 2916 -5013 2970 -5004
rect 2916 -5067 2970 -5058
rect 2916 -5103 2925 -5067
rect 2961 -5103 2970 -5067
rect 2916 -5112 2970 -5103
rect 3519 -5130 3564 -5121
rect 2916 -5139 2970 -5130
rect 2916 -5175 2925 -5139
rect 2961 -5175 2970 -5139
rect 2916 -5184 2970 -5175
rect 3519 -5148 3528 -5130
rect 3555 -5148 3564 -5130
rect 3582 -5148 3600 -5121
rect 3627 -5148 3636 -5121
rect 2916 -5256 2970 -5247
rect 2916 -5292 2925 -5256
rect 2961 -5292 2970 -5256
rect 2916 -5310 2970 -5292
rect 2916 -5337 2970 -5328
rect 2916 -5373 2925 -5337
rect 2961 -5373 2970 -5337
rect 2916 -5382 2970 -5373
rect 2916 -5418 2970 -5409
rect 2916 -5454 2925 -5418
rect 2961 -5454 2970 -5418
rect 2916 -5472 2970 -5454
rect 6624 -5193 6669 -5184
rect 6624 -5211 6633 -5193
rect 6660 -5211 6669 -5193
rect 6687 -5211 6705 -5184
rect 6732 -5211 6741 -5184
rect 6174 -5247 6210 -5238
rect 6174 -5265 6183 -5247
rect 6201 -5265 6210 -5247
rect 6228 -5265 6372 -5238
rect 6390 -5256 6399 -5238
rect 6417 -5256 6426 -5238
rect 6390 -5265 6426 -5256
rect 4824 -5301 4833 -5274
rect 4860 -5301 4869 -5274
rect 4887 -5301 4995 -5274
rect 5013 -5301 5139 -5274
rect 5157 -5301 5265 -5274
rect 5283 -5301 5400 -5274
rect 5418 -5301 5454 -5274
rect 5481 -5301 5553 -5274
rect 5607 -5301 5625 -5274
rect 5652 -5301 5661 -5274
rect 5679 -5301 5688 -5274
rect 5715 -5301 5724 -5274
rect 2916 -5499 2970 -5490
rect 2916 -5535 2925 -5499
rect 2961 -5535 2970 -5499
rect 2916 -5544 2970 -5535
rect 2916 -5913 2970 -5904
rect 2916 -5949 2925 -5913
rect 2961 -5949 2970 -5913
rect 2916 -5958 2970 -5949
rect 2916 -5985 2970 -5976
rect 2916 -6021 2925 -5985
rect 2961 -6021 2970 -5985
rect 2916 -6030 2970 -6021
rect 2916 -6084 2970 -6075
rect 2916 -6120 2925 -6084
rect 2961 -6120 2970 -6084
rect 2916 -6129 2970 -6120
rect 3519 -6147 3564 -6138
rect 2916 -6156 2970 -6147
rect 2916 -6192 2925 -6156
rect 2961 -6192 2970 -6156
rect 2916 -6201 2970 -6192
rect 3519 -6165 3528 -6147
rect 3555 -6165 3564 -6147
rect 3582 -6165 3600 -6138
rect 3627 -6165 3636 -6138
rect 2916 -6273 2970 -6264
rect 2916 -6309 2925 -6273
rect 2961 -6309 2970 -6273
rect 2916 -6327 2970 -6309
rect 2916 -6354 2970 -6345
rect 2916 -6390 2925 -6354
rect 2961 -6390 2970 -6354
rect 2916 -6399 2970 -6390
rect 2916 -6435 2970 -6426
rect 2916 -6471 2925 -6435
rect 2961 -6471 2970 -6435
rect 2916 -6489 2970 -6471
rect 2916 -6516 2970 -6507
rect 2916 -6552 2925 -6516
rect 2961 -6552 2970 -6516
rect 2916 -6561 2970 -6552
rect 2916 -7209 2970 -7200
rect 2916 -7245 2925 -7209
rect 2961 -7245 2970 -7209
rect 2916 -7254 2970 -7245
rect 2916 -7281 2970 -7272
rect 2916 -7317 2925 -7281
rect 2961 -7317 2970 -7281
rect 2916 -7326 2970 -7317
rect 2916 -7380 2970 -7371
rect 2916 -7416 2925 -7380
rect 2961 -7416 2970 -7380
rect 2916 -7425 2970 -7416
rect 3519 -7443 3564 -7434
rect 2916 -7452 2970 -7443
rect 2916 -7488 2925 -7452
rect 2961 -7488 2970 -7452
rect 2916 -7497 2970 -7488
rect 3519 -7461 3528 -7443
rect 3555 -7461 3564 -7443
rect 3582 -7461 3600 -7434
rect 3627 -7461 3636 -7434
rect 2916 -7569 2970 -7560
rect 2916 -7605 2925 -7569
rect 2961 -7605 2970 -7569
rect 2916 -7623 2970 -7605
rect 2916 -7650 2970 -7641
rect 2916 -7686 2925 -7650
rect 2961 -7686 2970 -7650
rect 2916 -7695 2970 -7686
rect 2916 -7731 2970 -7722
rect 2916 -7767 2925 -7731
rect 2961 -7767 2970 -7731
rect 2916 -7785 2970 -7767
rect 2916 -7812 2970 -7803
rect 2916 -7848 2925 -7812
rect 2961 -7848 2970 -7812
rect 2916 -7857 2970 -7848
<< pdiffusion >>
rect 3168 5175 3231 5184
rect 3168 5139 3177 5175
rect 3213 5139 3231 5175
rect 3168 5130 3231 5139
rect 3168 5103 3231 5112
rect 3168 5067 3177 5103
rect 3213 5067 3231 5103
rect 3168 5058 3231 5067
rect 3168 5004 3231 5013
rect 3168 4968 3177 5004
rect 3213 4968 3231 5004
rect 3168 4959 3231 4968
rect 3519 5049 3528 5076
rect 3555 5049 3564 5076
rect 3519 5022 3564 5049
rect 3582 5067 3636 5076
rect 3582 5040 3600 5067
rect 3627 5040 3636 5067
rect 3582 5022 3636 5040
rect 3168 4932 3231 4941
rect 3168 4896 3177 4932
rect 3213 4896 3231 4932
rect 3168 4887 3231 4896
rect 3168 4815 3231 4824
rect 3168 4779 3177 4815
rect 3213 4779 3231 4815
rect 3168 4761 3231 4779
rect 3168 4734 3231 4743
rect 3168 4698 3177 4734
rect 3213 4698 3231 4734
rect 3168 4689 3231 4698
rect 3168 4653 3231 4662
rect 3168 4617 3177 4653
rect 3213 4617 3231 4653
rect 3168 4599 3231 4617
rect 3168 4572 3231 4581
rect 3168 4536 3177 4572
rect 3213 4536 3231 4572
rect 3168 4527 3231 4536
rect 4725 4779 4734 4806
rect 4761 4779 4770 4806
rect 3888 4743 3897 4770
rect 3924 4743 3933 4770
rect 3888 4716 3933 4743
rect 3951 4761 4005 4770
rect 3951 4734 3969 4761
rect 3996 4734 4005 4761
rect 3951 4716 4005 4734
rect 4275 4761 4311 4770
rect 4275 4743 4284 4761
rect 4302 4743 4311 4761
rect 4275 4725 4311 4743
rect 4329 4752 4392 4770
rect 4329 4734 4338 4752
rect 4356 4734 4392 4752
rect 4329 4725 4392 4734
rect 4428 4761 4473 4770
rect 4428 4743 4437 4761
rect 4455 4743 4473 4761
rect 4428 4725 4473 4743
rect 4491 4761 4527 4770
rect 4491 4743 4500 4761
rect 4518 4743 4527 4761
rect 4725 4752 4770 4779
rect 4788 4797 4842 4806
rect 4788 4770 4806 4797
rect 4833 4770 4842 4797
rect 4788 4752 4842 4770
rect 4491 4725 4527 4743
rect 3168 4230 3231 4239
rect 3168 4194 3177 4230
rect 3213 4194 3231 4230
rect 3168 4185 3231 4194
rect 3168 4158 3231 4167
rect 3168 4122 3177 4158
rect 3213 4122 3231 4158
rect 3168 4113 3231 4122
rect 3168 4059 3231 4068
rect 3168 4023 3177 4059
rect 3213 4023 3231 4059
rect 3168 4014 3231 4023
rect 3519 4104 3528 4131
rect 3555 4104 3564 4131
rect 3519 4077 3564 4104
rect 3582 4122 3636 4131
rect 3582 4095 3600 4122
rect 3627 4095 3636 4122
rect 3582 4077 3636 4095
rect 3168 3987 3231 3996
rect 3168 3951 3177 3987
rect 3213 3951 3231 3987
rect 4653 3969 4662 3996
rect 4689 3969 4698 3996
rect 3168 3942 3231 3951
rect 3168 3870 3231 3879
rect 3168 3834 3177 3870
rect 3213 3834 3231 3870
rect 3168 3816 3231 3834
rect 3168 3789 3231 3798
rect 3168 3753 3177 3789
rect 3213 3753 3231 3789
rect 3870 3933 3879 3960
rect 3906 3933 3915 3960
rect 3870 3906 3915 3933
rect 3933 3951 3987 3960
rect 3933 3924 3951 3951
rect 3978 3924 3987 3951
rect 3933 3906 3987 3924
rect 4203 3951 4239 3960
rect 4203 3933 4212 3951
rect 4230 3933 4239 3951
rect 4203 3915 4239 3933
rect 4257 3942 4320 3960
rect 4257 3924 4266 3942
rect 4284 3924 4320 3942
rect 4257 3915 4320 3924
rect 4356 3951 4401 3960
rect 4356 3933 4365 3951
rect 4383 3933 4401 3951
rect 4356 3915 4401 3933
rect 4419 3951 4455 3960
rect 4419 3933 4428 3951
rect 4446 3933 4455 3951
rect 4653 3942 4698 3969
rect 4716 3987 4770 3996
rect 4716 3960 4734 3987
rect 4761 3960 4770 3987
rect 4716 3942 4770 3960
rect 5031 3951 5067 3960
rect 4419 3915 4455 3933
rect 5031 3933 5040 3951
rect 5058 3933 5067 3951
rect 5031 3915 5067 3933
rect 5085 3942 5148 3960
rect 5085 3924 5094 3942
rect 5112 3924 5148 3942
rect 5085 3915 5148 3924
rect 5481 3969 5490 3996
rect 5517 3969 5526 3996
rect 5184 3951 5229 3960
rect 5184 3933 5193 3951
rect 5211 3933 5229 3951
rect 5184 3915 5229 3933
rect 5247 3951 5283 3960
rect 5247 3933 5256 3951
rect 5274 3933 5283 3951
rect 5481 3942 5526 3969
rect 5544 3987 5598 3996
rect 5544 3960 5562 3987
rect 5589 3960 5598 3987
rect 5544 3942 5598 3960
rect 5904 3942 5949 3951
rect 5247 3915 5283 3933
rect 5904 3924 5913 3942
rect 5931 3924 5949 3942
rect 5904 3906 5949 3924
rect 5967 3906 6003 3951
rect 6021 3906 6039 3951
rect 6057 3906 6129 3951
rect 6147 3906 6219 3951
rect 6237 3933 6264 3951
rect 6237 3915 6246 3933
rect 6237 3906 6264 3915
rect 6309 3942 6345 3951
rect 6309 3924 6318 3942
rect 6336 3924 6345 3942
rect 6309 3906 6345 3924
rect 6363 3933 6399 3951
rect 6363 3915 6372 3933
rect 6390 3915 6399 3933
rect 6363 3906 6399 3915
rect 3168 3744 3231 3753
rect 3168 3708 3231 3717
rect 3168 3672 3177 3708
rect 3213 3672 3231 3708
rect 3168 3654 3231 3672
rect 3168 3627 3231 3636
rect 3168 3591 3177 3627
rect 3213 3591 3231 3627
rect 3168 3582 3231 3591
rect 3168 3213 3231 3222
rect 3168 3177 3177 3213
rect 3213 3177 3231 3213
rect 3168 3168 3231 3177
rect 3168 3141 3231 3150
rect 3168 3105 3177 3141
rect 3213 3105 3231 3141
rect 3168 3096 3231 3105
rect 3168 3042 3231 3051
rect 3168 3006 3177 3042
rect 3213 3006 3231 3042
rect 3168 2997 3231 3006
rect 4356 3177 4401 3186
rect 4356 3150 4365 3177
rect 4392 3150 4401 3177
rect 4356 3132 4401 3150
rect 4419 3168 4464 3186
rect 4419 3141 4428 3168
rect 4455 3141 4464 3168
rect 4419 3132 4464 3141
rect 4482 3177 4527 3186
rect 4482 3150 4491 3177
rect 4518 3150 4527 3177
rect 4482 3132 4527 3150
rect 4545 3168 4599 3186
rect 4545 3141 4554 3168
rect 4581 3141 4599 3168
rect 4545 3132 4599 3141
rect 4617 3177 4671 3186
rect 4617 3150 4635 3177
rect 4662 3150 4671 3177
rect 4617 3132 4671 3150
rect 4689 3168 4734 3186
rect 4689 3141 4698 3168
rect 4725 3141 4734 3168
rect 4689 3132 4734 3141
rect 4752 3177 4797 3186
rect 4752 3150 4761 3177
rect 4788 3150 4797 3177
rect 4752 3132 4797 3150
rect 4815 3168 4860 3186
rect 4815 3141 4824 3168
rect 4851 3141 4860 3168
rect 4815 3132 4860 3141
rect 4878 3177 4932 3186
rect 4878 3150 4887 3177
rect 4914 3150 4932 3177
rect 4878 3132 4932 3150
rect 4950 3168 5085 3186
rect 4950 3141 4959 3168
rect 4986 3141 5085 3168
rect 4950 3132 5085 3141
rect 5139 3159 5157 3186
rect 5184 3159 5193 3186
rect 5139 3132 5193 3159
rect 5211 3168 5256 3186
rect 5211 3141 5220 3168
rect 5247 3141 5256 3168
rect 5211 3132 5256 3141
rect 3519 3087 3528 3114
rect 3555 3087 3564 3114
rect 3519 3060 3564 3087
rect 3582 3105 3636 3114
rect 3582 3078 3600 3105
rect 3627 3078 3636 3105
rect 3582 3060 3636 3078
rect 3852 3087 3861 3114
rect 3888 3087 3897 3114
rect 3852 3060 3897 3087
rect 3915 3105 3969 3114
rect 3915 3078 3933 3105
rect 3960 3078 3969 3105
rect 3915 3060 3969 3078
rect 3168 2970 3231 2979
rect 3168 2934 3177 2970
rect 3213 2934 3231 2970
rect 3168 2925 3231 2934
rect 3168 2853 3231 2862
rect 3168 2817 3177 2853
rect 3213 2817 3231 2853
rect 3168 2799 3231 2817
rect 3168 2772 3231 2781
rect 3168 2736 3177 2772
rect 3213 2736 3231 2772
rect 3168 2727 3231 2736
rect 3168 2691 3231 2700
rect 3168 2655 3177 2691
rect 3213 2655 3231 2691
rect 3168 2637 3231 2655
rect 3168 2610 3231 2619
rect 3168 2574 3177 2610
rect 3213 2574 3231 2610
rect 3168 2565 3231 2574
rect 3168 1917 3231 1926
rect 3168 1881 3177 1917
rect 3213 1881 3231 1917
rect 3168 1872 3231 1881
rect 3168 1845 3231 1854
rect 3168 1809 3177 1845
rect 3213 1809 3231 1845
rect 3168 1800 3231 1809
rect 3168 1746 3231 1755
rect 3168 1710 3177 1746
rect 3213 1710 3231 1746
rect 3168 1701 3231 1710
rect 4203 1881 4248 1890
rect 4203 1854 4212 1881
rect 4239 1854 4248 1881
rect 4203 1836 4248 1854
rect 4266 1872 4311 1890
rect 4266 1845 4275 1872
rect 4302 1845 4311 1872
rect 4266 1836 4311 1845
rect 4329 1881 4374 1890
rect 4329 1854 4338 1881
rect 4365 1854 4374 1881
rect 4329 1836 4374 1854
rect 4392 1872 4446 1890
rect 4392 1845 4401 1872
rect 4428 1845 4446 1872
rect 4392 1836 4446 1845
rect 4464 1881 4518 1890
rect 4464 1854 4482 1881
rect 4509 1854 4518 1881
rect 4464 1836 4518 1854
rect 4536 1872 4581 1890
rect 4536 1845 4545 1872
rect 4572 1845 4581 1872
rect 4536 1836 4581 1845
rect 4599 1881 4644 1890
rect 4599 1854 4608 1881
rect 4635 1854 4644 1881
rect 4599 1836 4644 1854
rect 4662 1872 4707 1890
rect 4662 1845 4671 1872
rect 4698 1845 4707 1872
rect 4662 1836 4707 1845
rect 4725 1881 4779 1890
rect 4725 1854 4734 1881
rect 4761 1854 4779 1881
rect 4725 1836 4779 1854
rect 4797 1872 4932 1890
rect 4797 1845 4806 1872
rect 4833 1845 4932 1872
rect 4797 1836 4932 1845
rect 4986 1863 5004 1890
rect 5031 1863 5040 1890
rect 4986 1836 5040 1863
rect 5058 1872 5103 1890
rect 5058 1845 5067 1872
rect 5094 1845 5103 1872
rect 5058 1836 5103 1845
rect 3519 1791 3528 1818
rect 3555 1791 3564 1818
rect 3519 1764 3564 1791
rect 3582 1809 3636 1818
rect 3582 1782 3600 1809
rect 3627 1782 3636 1809
rect 3582 1764 3636 1782
rect 3798 1791 3807 1818
rect 3834 1791 3843 1818
rect 3798 1764 3843 1791
rect 3861 1809 3915 1818
rect 3861 1782 3879 1809
rect 3906 1782 3915 1809
rect 3861 1764 3915 1782
rect 3168 1674 3231 1683
rect 3168 1638 3177 1674
rect 3213 1638 3231 1674
rect 3168 1629 3231 1638
rect 3168 1557 3231 1566
rect 3168 1521 3177 1557
rect 3213 1521 3231 1557
rect 3168 1503 3231 1521
rect 3168 1476 3231 1485
rect 3168 1440 3177 1476
rect 3213 1440 3231 1476
rect 3168 1431 3231 1440
rect 3168 1395 3231 1404
rect 3168 1359 3177 1395
rect 3213 1359 3231 1395
rect 3168 1341 3231 1359
rect 3168 1314 3231 1323
rect 3168 1278 3177 1314
rect 3213 1278 3231 1314
rect 3168 1269 3231 1278
rect 3168 846 3231 855
rect 3168 810 3177 846
rect 3213 810 3231 846
rect 3168 801 3231 810
rect 3168 774 3231 783
rect 3168 738 3177 774
rect 3213 738 3231 774
rect 3168 729 3231 738
rect 3168 675 3231 684
rect 3168 639 3177 675
rect 3213 639 3231 675
rect 3168 630 3231 639
rect 3519 720 3528 747
rect 3555 720 3564 747
rect 3519 693 3564 720
rect 3582 738 3636 747
rect 3582 711 3600 738
rect 3627 711 3636 738
rect 3582 693 3636 711
rect 3168 603 3231 612
rect 3168 567 3177 603
rect 3213 567 3231 603
rect 3168 558 3231 567
rect 3168 486 3231 495
rect 3168 450 3177 486
rect 3213 450 3231 486
rect 3168 432 3231 450
rect 3168 405 3231 414
rect 3168 369 3177 405
rect 3213 369 3231 405
rect 3168 360 3231 369
rect 3168 324 3231 333
rect 3168 288 3177 324
rect 3213 288 3231 324
rect 3168 270 3231 288
rect 3168 243 3231 252
rect 3168 207 3177 243
rect 3213 207 3231 243
rect 3168 198 3231 207
rect 4725 450 4734 477
rect 4761 450 4770 477
rect 3888 414 3897 441
rect 3924 414 3933 441
rect 3888 387 3933 414
rect 3951 432 4005 441
rect 3951 405 3969 432
rect 3996 405 4005 432
rect 3951 387 4005 405
rect 4275 432 4311 441
rect 4275 414 4284 432
rect 4302 414 4311 432
rect 4275 396 4311 414
rect 4329 423 4392 441
rect 4329 405 4338 423
rect 4356 405 4392 423
rect 4329 396 4392 405
rect 4428 432 4473 441
rect 4428 414 4437 432
rect 4455 414 4473 432
rect 4428 396 4473 414
rect 4491 432 4527 441
rect 4491 414 4500 432
rect 4518 414 4527 432
rect 4725 423 4770 450
rect 4788 468 4842 477
rect 4788 441 4806 468
rect 4833 441 4842 468
rect 4788 423 4842 441
rect 4491 396 4527 414
rect 3168 -99 3231 -90
rect 3168 -135 3177 -99
rect 3213 -135 3231 -99
rect 3168 -144 3231 -135
rect 3168 -171 3231 -162
rect 3168 -207 3177 -171
rect 3213 -207 3231 -171
rect 3168 -216 3231 -207
rect 3168 -270 3231 -261
rect 3168 -306 3177 -270
rect 3213 -306 3231 -270
rect 3168 -315 3231 -306
rect 3519 -225 3528 -198
rect 3555 -225 3564 -198
rect 3519 -252 3564 -225
rect 3582 -207 3636 -198
rect 3582 -234 3600 -207
rect 3627 -234 3636 -207
rect 3582 -252 3636 -234
rect 3168 -342 3231 -333
rect 3168 -378 3177 -342
rect 3213 -378 3231 -342
rect 4653 -360 4662 -333
rect 4689 -360 4698 -333
rect 3168 -387 3231 -378
rect 3168 -459 3231 -450
rect 3168 -495 3177 -459
rect 3213 -495 3231 -459
rect 3168 -513 3231 -495
rect 3168 -540 3231 -531
rect 3168 -576 3177 -540
rect 3213 -576 3231 -540
rect 3870 -396 3879 -369
rect 3906 -396 3915 -369
rect 3870 -423 3915 -396
rect 3933 -378 3987 -369
rect 3933 -405 3951 -378
rect 3978 -405 3987 -378
rect 3933 -423 3987 -405
rect 4203 -378 4239 -369
rect 4203 -396 4212 -378
rect 4230 -396 4239 -378
rect 4203 -414 4239 -396
rect 4257 -387 4320 -369
rect 4257 -405 4266 -387
rect 4284 -405 4320 -387
rect 4257 -414 4320 -405
rect 4356 -378 4401 -369
rect 4356 -396 4365 -378
rect 4383 -396 4401 -378
rect 4356 -414 4401 -396
rect 4419 -378 4455 -369
rect 4419 -396 4428 -378
rect 4446 -396 4455 -378
rect 4653 -387 4698 -360
rect 4716 -342 4770 -333
rect 4716 -369 4734 -342
rect 4761 -369 4770 -342
rect 4716 -387 4770 -369
rect 5031 -378 5067 -369
rect 4419 -414 4455 -396
rect 5031 -396 5040 -378
rect 5058 -396 5067 -378
rect 5031 -414 5067 -396
rect 5085 -387 5148 -369
rect 5085 -405 5094 -387
rect 5112 -405 5148 -387
rect 5085 -414 5148 -405
rect 5481 -360 5490 -333
rect 5517 -360 5526 -333
rect 5184 -378 5229 -369
rect 5184 -396 5193 -378
rect 5211 -396 5229 -378
rect 5184 -414 5229 -396
rect 5247 -378 5283 -369
rect 5247 -396 5256 -378
rect 5274 -396 5283 -378
rect 5481 -387 5526 -360
rect 5544 -342 5598 -333
rect 5544 -369 5562 -342
rect 5589 -369 5598 -342
rect 5544 -387 5598 -369
rect 5904 -387 5949 -378
rect 5247 -414 5283 -396
rect 5904 -405 5913 -387
rect 5931 -405 5949 -387
rect 5904 -423 5949 -405
rect 5967 -423 6003 -378
rect 6021 -423 6039 -378
rect 6057 -423 6129 -378
rect 6147 -423 6219 -378
rect 6237 -396 6264 -378
rect 6237 -414 6246 -396
rect 6237 -423 6264 -414
rect 6309 -387 6345 -378
rect 6309 -405 6318 -387
rect 6336 -405 6345 -387
rect 6309 -423 6345 -405
rect 6363 -396 6399 -378
rect 6363 -414 6372 -396
rect 6390 -414 6399 -396
rect 6363 -423 6399 -414
rect 3168 -585 3231 -576
rect 3168 -621 3231 -612
rect 3168 -657 3177 -621
rect 3213 -657 3231 -621
rect 3168 -675 3231 -657
rect 3168 -702 3231 -693
rect 3168 -738 3177 -702
rect 3213 -738 3231 -702
rect 3168 -747 3231 -738
rect 3168 -1116 3231 -1107
rect 3168 -1152 3177 -1116
rect 3213 -1152 3231 -1116
rect 3168 -1161 3231 -1152
rect 3168 -1188 3231 -1179
rect 3168 -1224 3177 -1188
rect 3213 -1224 3231 -1188
rect 3168 -1233 3231 -1224
rect 3168 -1287 3231 -1278
rect 3168 -1323 3177 -1287
rect 3213 -1323 3231 -1287
rect 3168 -1332 3231 -1323
rect 4356 -1152 4401 -1143
rect 4356 -1179 4365 -1152
rect 4392 -1179 4401 -1152
rect 4356 -1197 4401 -1179
rect 4419 -1161 4464 -1143
rect 4419 -1188 4428 -1161
rect 4455 -1188 4464 -1161
rect 4419 -1197 4464 -1188
rect 4482 -1152 4527 -1143
rect 4482 -1179 4491 -1152
rect 4518 -1179 4527 -1152
rect 4482 -1197 4527 -1179
rect 4545 -1161 4599 -1143
rect 4545 -1188 4554 -1161
rect 4581 -1188 4599 -1161
rect 4545 -1197 4599 -1188
rect 4617 -1152 4671 -1143
rect 4617 -1179 4635 -1152
rect 4662 -1179 4671 -1152
rect 4617 -1197 4671 -1179
rect 4689 -1161 4734 -1143
rect 4689 -1188 4698 -1161
rect 4725 -1188 4734 -1161
rect 4689 -1197 4734 -1188
rect 4752 -1152 4797 -1143
rect 4752 -1179 4761 -1152
rect 4788 -1179 4797 -1152
rect 4752 -1197 4797 -1179
rect 4815 -1161 4860 -1143
rect 4815 -1188 4824 -1161
rect 4851 -1188 4860 -1161
rect 4815 -1197 4860 -1188
rect 4878 -1152 4932 -1143
rect 4878 -1179 4887 -1152
rect 4914 -1179 4932 -1152
rect 4878 -1197 4932 -1179
rect 4950 -1161 5085 -1143
rect 4950 -1188 4959 -1161
rect 4986 -1188 5085 -1161
rect 4950 -1197 5085 -1188
rect 5139 -1170 5157 -1143
rect 5184 -1170 5193 -1143
rect 5139 -1197 5193 -1170
rect 5211 -1161 5256 -1143
rect 5211 -1188 5220 -1161
rect 5247 -1188 5256 -1161
rect 5211 -1197 5256 -1188
rect 3519 -1242 3528 -1215
rect 3555 -1242 3564 -1215
rect 3519 -1269 3564 -1242
rect 3582 -1224 3636 -1215
rect 3582 -1251 3600 -1224
rect 3627 -1251 3636 -1224
rect 3582 -1269 3636 -1251
rect 3852 -1242 3861 -1215
rect 3888 -1242 3897 -1215
rect 3852 -1269 3897 -1242
rect 3915 -1224 3969 -1215
rect 3915 -1251 3933 -1224
rect 3960 -1251 3969 -1224
rect 3915 -1269 3969 -1251
rect 3168 -1359 3231 -1350
rect 3168 -1395 3177 -1359
rect 3213 -1395 3231 -1359
rect 3168 -1404 3231 -1395
rect 3168 -1476 3231 -1467
rect 3168 -1512 3177 -1476
rect 3213 -1512 3231 -1476
rect 3168 -1530 3231 -1512
rect 3168 -1557 3231 -1548
rect 3168 -1593 3177 -1557
rect 3213 -1593 3231 -1557
rect 3168 -1602 3231 -1593
rect 3168 -1638 3231 -1629
rect 3168 -1674 3177 -1638
rect 3213 -1674 3231 -1638
rect 3168 -1692 3231 -1674
rect 3168 -1719 3231 -1710
rect 3168 -1755 3177 -1719
rect 3213 -1755 3231 -1719
rect 3168 -1764 3231 -1755
rect 3168 -2412 3231 -2403
rect 3168 -2448 3177 -2412
rect 3213 -2448 3231 -2412
rect 3168 -2457 3231 -2448
rect 3168 -2484 3231 -2475
rect 3168 -2520 3177 -2484
rect 3213 -2520 3231 -2484
rect 3168 -2529 3231 -2520
rect 3168 -2583 3231 -2574
rect 3168 -2619 3177 -2583
rect 3213 -2619 3231 -2583
rect 3168 -2628 3231 -2619
rect 3519 -2538 3528 -2511
rect 3555 -2538 3564 -2511
rect 3519 -2565 3564 -2538
rect 3582 -2520 3636 -2511
rect 3582 -2547 3600 -2520
rect 3627 -2547 3636 -2520
rect 3582 -2565 3636 -2547
rect 3168 -2655 3231 -2646
rect 3168 -2691 3177 -2655
rect 3213 -2691 3231 -2655
rect 3168 -2700 3231 -2691
rect 3168 -2772 3231 -2763
rect 3168 -2808 3177 -2772
rect 3213 -2808 3231 -2772
rect 3168 -2826 3231 -2808
rect 3168 -2853 3231 -2844
rect 3168 -2889 3177 -2853
rect 3213 -2889 3231 -2853
rect 3168 -2898 3231 -2889
rect 3168 -2934 3231 -2925
rect 3168 -2970 3177 -2934
rect 3213 -2970 3231 -2934
rect 3168 -2988 3231 -2970
rect 3168 -3015 3231 -3006
rect 3168 -3051 3177 -3015
rect 3213 -3051 3231 -3015
rect 3168 -3060 3231 -3051
rect 3168 -3951 3231 -3942
rect 3168 -3987 3177 -3951
rect 3213 -3987 3231 -3951
rect 3168 -3996 3231 -3987
rect 3168 -4023 3231 -4014
rect 3168 -4059 3177 -4023
rect 3213 -4059 3231 -4023
rect 3168 -4068 3231 -4059
rect 3168 -4122 3231 -4113
rect 3168 -4158 3177 -4122
rect 3213 -4158 3231 -4122
rect 3168 -4167 3231 -4158
rect 4203 -2448 4248 -2439
rect 4203 -2475 4212 -2448
rect 4239 -2475 4248 -2448
rect 4203 -2493 4248 -2475
rect 4266 -2457 4311 -2439
rect 4266 -2484 4275 -2457
rect 4302 -2484 4311 -2457
rect 4266 -2493 4311 -2484
rect 4329 -2448 4374 -2439
rect 4329 -2475 4338 -2448
rect 4365 -2475 4374 -2448
rect 4329 -2493 4374 -2475
rect 4392 -2457 4446 -2439
rect 4392 -2484 4401 -2457
rect 4428 -2484 4446 -2457
rect 4392 -2493 4446 -2484
rect 4464 -2448 4518 -2439
rect 4464 -2475 4482 -2448
rect 4509 -2475 4518 -2448
rect 4464 -2493 4518 -2475
rect 4536 -2457 4581 -2439
rect 4536 -2484 4545 -2457
rect 4572 -2484 4581 -2457
rect 4536 -2493 4581 -2484
rect 4599 -2448 4644 -2439
rect 4599 -2475 4608 -2448
rect 4635 -2475 4644 -2448
rect 4599 -2493 4644 -2475
rect 4662 -2457 4707 -2439
rect 4662 -2484 4671 -2457
rect 4698 -2484 4707 -2457
rect 4662 -2493 4707 -2484
rect 4725 -2448 4779 -2439
rect 4725 -2475 4734 -2448
rect 4761 -2475 4779 -2448
rect 4725 -2493 4779 -2475
rect 4797 -2457 4932 -2439
rect 4797 -2484 4806 -2457
rect 4833 -2484 4932 -2457
rect 4797 -2493 4932 -2484
rect 4986 -2466 5004 -2439
rect 5031 -2466 5040 -2439
rect 4986 -2493 5040 -2466
rect 5058 -2457 5103 -2439
rect 5058 -2484 5067 -2457
rect 5094 -2484 5103 -2457
rect 5058 -2493 5103 -2484
rect 3798 -2538 3807 -2511
rect 3834 -2538 3843 -2511
rect 3798 -2565 3843 -2538
rect 3861 -2520 3915 -2511
rect 3861 -2547 3879 -2520
rect 3906 -2547 3915 -2520
rect 3861 -2565 3915 -2547
rect 3519 -4077 3528 -4050
rect 3555 -4077 3564 -4050
rect 3519 -4104 3564 -4077
rect 3582 -4059 3636 -4050
rect 3582 -4086 3600 -4059
rect 3627 -4086 3636 -4059
rect 3582 -4104 3636 -4086
rect 3168 -4194 3231 -4185
rect 3168 -4230 3177 -4194
rect 3213 -4230 3231 -4194
rect 3168 -4239 3231 -4230
rect 3168 -4311 3231 -4302
rect 3168 -4347 3177 -4311
rect 3213 -4347 3231 -4311
rect 3168 -4365 3231 -4347
rect 3168 -4392 3231 -4383
rect 3168 -4428 3177 -4392
rect 3213 -4428 3231 -4392
rect 3168 -4437 3231 -4428
rect 3168 -4473 3231 -4464
rect 3168 -4509 3177 -4473
rect 3213 -4509 3231 -4473
rect 3168 -4527 3231 -4509
rect 3168 -4554 3231 -4545
rect 3168 -4590 3177 -4554
rect 3213 -4590 3231 -4554
rect 3168 -4599 3231 -4590
rect 3168 -4896 3231 -4887
rect 3168 -4932 3177 -4896
rect 3213 -4932 3231 -4896
rect 3168 -4941 3231 -4932
rect 3168 -4968 3231 -4959
rect 3168 -5004 3177 -4968
rect 3213 -5004 3231 -4968
rect 3168 -5013 3231 -5004
rect 3168 -5067 3231 -5058
rect 3168 -5103 3177 -5067
rect 3213 -5103 3231 -5067
rect 3168 -5112 3231 -5103
rect 3519 -5022 3528 -4995
rect 3555 -5022 3564 -4995
rect 3519 -5049 3564 -5022
rect 3582 -5004 3636 -4995
rect 3582 -5031 3600 -5004
rect 3627 -5031 3636 -5004
rect 3582 -5049 3636 -5031
rect 3168 -5139 3231 -5130
rect 3168 -5175 3177 -5139
rect 3213 -5175 3231 -5139
rect 3168 -5184 3231 -5175
rect 3168 -5256 3231 -5247
rect 3168 -5292 3177 -5256
rect 3213 -5292 3231 -5256
rect 3168 -5310 3231 -5292
rect 3168 -5337 3231 -5328
rect 3168 -5373 3177 -5337
rect 3213 -5373 3231 -5337
rect 3168 -5382 3231 -5373
rect 3168 -5418 3231 -5409
rect 3168 -5454 3177 -5418
rect 3213 -5454 3231 -5418
rect 6624 -5085 6633 -5058
rect 6660 -5085 6669 -5058
rect 4824 -5103 4869 -5094
rect 4824 -5130 4833 -5103
rect 4860 -5130 4869 -5103
rect 4824 -5148 4869 -5130
rect 4887 -5112 4932 -5094
rect 4887 -5139 4896 -5112
rect 4923 -5139 4932 -5112
rect 4887 -5148 4932 -5139
rect 4950 -5103 4995 -5094
rect 4950 -5130 4959 -5103
rect 4986 -5130 4995 -5103
rect 4950 -5148 4995 -5130
rect 5013 -5112 5067 -5094
rect 5013 -5139 5022 -5112
rect 5049 -5139 5067 -5112
rect 5013 -5148 5067 -5139
rect 5085 -5103 5139 -5094
rect 5085 -5130 5103 -5103
rect 5130 -5130 5139 -5103
rect 5085 -5148 5139 -5130
rect 5157 -5112 5202 -5094
rect 5157 -5139 5166 -5112
rect 5193 -5139 5202 -5112
rect 5157 -5148 5202 -5139
rect 5220 -5103 5265 -5094
rect 5220 -5130 5229 -5103
rect 5256 -5130 5265 -5103
rect 5220 -5148 5265 -5130
rect 5283 -5112 5328 -5094
rect 5283 -5139 5292 -5112
rect 5319 -5139 5328 -5112
rect 5283 -5148 5328 -5139
rect 5346 -5103 5400 -5094
rect 5346 -5130 5355 -5103
rect 5382 -5130 5400 -5103
rect 5346 -5148 5400 -5130
rect 5418 -5112 5553 -5094
rect 5418 -5139 5427 -5112
rect 5454 -5139 5553 -5112
rect 5418 -5148 5553 -5139
rect 5607 -5121 5625 -5094
rect 5652 -5121 5661 -5094
rect 5607 -5148 5661 -5121
rect 5679 -5112 5724 -5094
rect 5679 -5139 5688 -5112
rect 5715 -5139 5724 -5112
rect 6174 -5103 6210 -5094
rect 6174 -5121 6183 -5103
rect 6201 -5121 6210 -5103
rect 6174 -5139 6210 -5121
rect 6228 -5112 6291 -5094
rect 6228 -5130 6237 -5112
rect 6255 -5130 6291 -5112
rect 6228 -5139 6291 -5130
rect 6327 -5103 6372 -5094
rect 6327 -5121 6336 -5103
rect 6354 -5121 6372 -5103
rect 6327 -5139 6372 -5121
rect 6390 -5103 6426 -5094
rect 6390 -5121 6399 -5103
rect 6417 -5121 6426 -5103
rect 6624 -5112 6669 -5085
rect 6687 -5067 6741 -5058
rect 6687 -5094 6705 -5067
rect 6732 -5094 6741 -5067
rect 6687 -5112 6741 -5094
rect 6390 -5139 6426 -5121
rect 5679 -5148 5724 -5139
rect 3168 -5472 3231 -5454
rect 3168 -5499 3231 -5490
rect 3168 -5535 3177 -5499
rect 3213 -5535 3231 -5499
rect 3168 -5544 3231 -5535
rect 3168 -5913 3231 -5904
rect 3168 -5949 3177 -5913
rect 3213 -5949 3231 -5913
rect 3168 -5958 3231 -5949
rect 3168 -5985 3231 -5976
rect 3168 -6021 3177 -5985
rect 3213 -6021 3231 -5985
rect 3168 -6030 3231 -6021
rect 3168 -6084 3231 -6075
rect 3168 -6120 3177 -6084
rect 3213 -6120 3231 -6084
rect 3168 -6129 3231 -6120
rect 3519 -6039 3528 -6012
rect 3555 -6039 3564 -6012
rect 3519 -6066 3564 -6039
rect 3582 -6021 3636 -6012
rect 3582 -6048 3600 -6021
rect 3627 -6048 3636 -6021
rect 3582 -6066 3636 -6048
rect 3168 -6156 3231 -6147
rect 3168 -6192 3177 -6156
rect 3213 -6192 3231 -6156
rect 3168 -6201 3231 -6192
rect 3168 -6273 3231 -6264
rect 3168 -6309 3177 -6273
rect 3213 -6309 3231 -6273
rect 3168 -6327 3231 -6309
rect 3168 -6354 3231 -6345
rect 3168 -6390 3177 -6354
rect 3213 -6390 3231 -6354
rect 3168 -6399 3231 -6390
rect 3168 -6435 3231 -6426
rect 3168 -6471 3177 -6435
rect 3213 -6471 3231 -6435
rect 3168 -6489 3231 -6471
rect 3168 -6516 3231 -6507
rect 3168 -6552 3177 -6516
rect 3213 -6552 3231 -6516
rect 3168 -6561 3231 -6552
rect 3168 -7209 3231 -7200
rect 3168 -7245 3177 -7209
rect 3213 -7245 3231 -7209
rect 3168 -7254 3231 -7245
rect 3168 -7281 3231 -7272
rect 3168 -7317 3177 -7281
rect 3213 -7317 3231 -7281
rect 3168 -7326 3231 -7317
rect 3168 -7380 3231 -7371
rect 3168 -7416 3177 -7380
rect 3213 -7416 3231 -7380
rect 3168 -7425 3231 -7416
rect 3519 -7335 3528 -7308
rect 3555 -7335 3564 -7308
rect 3519 -7362 3564 -7335
rect 3582 -7317 3636 -7308
rect 3582 -7344 3600 -7317
rect 3627 -7344 3636 -7317
rect 3582 -7362 3636 -7344
rect 3168 -7452 3231 -7443
rect 3168 -7488 3177 -7452
rect 3213 -7488 3231 -7452
rect 3168 -7497 3231 -7488
rect 3168 -7569 3231 -7560
rect 3168 -7605 3177 -7569
rect 3213 -7605 3231 -7569
rect 3168 -7623 3231 -7605
rect 3168 -7650 3231 -7641
rect 3168 -7686 3177 -7650
rect 3213 -7686 3231 -7650
rect 3168 -7695 3231 -7686
rect 3168 -7731 3231 -7722
rect 3168 -7767 3177 -7731
rect 3213 -7767 3231 -7731
rect 3168 -7785 3231 -7767
rect 3168 -7812 3231 -7803
rect 3168 -7848 3177 -7812
rect 3213 -7848 3231 -7812
rect 3168 -7857 3231 -7848
<< ndcontact >>
rect 2925 5139 2961 5175
rect 2925 5067 2961 5103
rect 2925 4968 2961 5004
rect 2925 4896 2961 4932
rect 3528 4914 3555 4941
rect 3600 4923 3627 4950
rect 2925 4779 2961 4815
rect 2925 4698 2961 4734
rect 2925 4617 2961 4653
rect 2925 4536 2961 4572
rect 3897 4608 3924 4635
rect 3969 4617 3996 4644
rect 4734 4644 4761 4671
rect 4806 4653 4833 4680
rect 4284 4599 4302 4617
rect 4500 4608 4518 4626
rect 2925 4194 2961 4230
rect 2925 4122 2961 4158
rect 2925 4023 2961 4059
rect 2925 3951 2961 3987
rect 3528 3969 3555 3996
rect 3600 3978 3627 4005
rect 2925 3834 2961 3870
rect 2925 3753 2961 3789
rect 3879 3798 3906 3825
rect 3951 3807 3978 3834
rect 4662 3834 4689 3861
rect 4734 3843 4761 3870
rect 5490 3834 5517 3861
rect 5562 3843 5589 3870
rect 4212 3789 4230 3807
rect 4428 3798 4446 3816
rect 5040 3789 5058 3807
rect 5256 3798 5274 3816
rect 5913 3798 5931 3816
rect 5976 3798 5994 3816
rect 6012 3798 6030 3816
rect 6066 3798 6084 3816
rect 6102 3798 6120 3816
rect 6156 3798 6174 3816
rect 6192 3798 6210 3816
rect 6246 3798 6264 3816
rect 6318 3798 6336 3816
rect 6372 3798 6390 3816
rect 2925 3672 2961 3708
rect 2925 3591 2961 3627
rect 2925 3177 2961 3213
rect 2925 3105 2961 3141
rect 2925 3006 2961 3042
rect 2925 2934 2961 2970
rect 3528 2952 3555 2979
rect 3600 2961 3627 2988
rect 3861 2952 3888 2979
rect 3933 2961 3960 2988
rect 4365 2979 4392 3006
rect 4986 2979 5013 3006
rect 5157 2979 5184 3006
rect 5220 2979 5247 3006
rect 2925 2817 2961 2853
rect 2925 2736 2961 2772
rect 2925 2655 2961 2691
rect 2925 2574 2961 2610
rect 2925 1881 2961 1917
rect 2925 1809 2961 1845
rect 2925 1710 2961 1746
rect 2925 1638 2961 1674
rect 3528 1656 3555 1683
rect 3600 1665 3627 1692
rect 3807 1656 3834 1683
rect 3879 1665 3906 1692
rect 4212 1683 4239 1710
rect 4833 1683 4860 1710
rect 5004 1683 5031 1710
rect 5067 1683 5094 1710
rect 2925 1521 2961 1557
rect 2925 1440 2961 1476
rect 2925 1359 2961 1395
rect 2925 1278 2961 1314
rect 2925 810 2961 846
rect 2925 738 2961 774
rect 2925 639 2961 675
rect 2925 567 2961 603
rect 3528 585 3555 612
rect 3600 594 3627 621
rect 2925 450 2961 486
rect 2925 369 2961 405
rect 2925 288 2961 324
rect 2925 207 2961 243
rect 3897 279 3924 306
rect 3969 288 3996 315
rect 4734 315 4761 342
rect 4806 324 4833 351
rect 4284 270 4302 288
rect 4500 279 4518 297
rect 2925 -135 2961 -99
rect 2925 -207 2961 -171
rect 2925 -306 2961 -270
rect 2925 -378 2961 -342
rect 3528 -360 3555 -333
rect 3600 -351 3627 -324
rect 2925 -495 2961 -459
rect 2925 -576 2961 -540
rect 3879 -531 3906 -504
rect 3951 -522 3978 -495
rect 4662 -495 4689 -468
rect 4734 -486 4761 -459
rect 5490 -495 5517 -468
rect 5562 -486 5589 -459
rect 4212 -540 4230 -522
rect 4428 -531 4446 -513
rect 5040 -540 5058 -522
rect 5256 -531 5274 -513
rect 5913 -531 5931 -513
rect 5976 -531 5994 -513
rect 6012 -531 6030 -513
rect 6066 -531 6084 -513
rect 6102 -531 6120 -513
rect 6156 -531 6174 -513
rect 6192 -531 6210 -513
rect 6246 -531 6264 -513
rect 6318 -531 6336 -513
rect 6372 -531 6390 -513
rect 2925 -657 2961 -621
rect 2925 -738 2961 -702
rect 2925 -1152 2961 -1116
rect 2925 -1224 2961 -1188
rect 2925 -1323 2961 -1287
rect 2925 -1395 2961 -1359
rect 3528 -1377 3555 -1350
rect 3600 -1368 3627 -1341
rect 3861 -1377 3888 -1350
rect 3933 -1368 3960 -1341
rect 4365 -1350 4392 -1323
rect 4986 -1350 5013 -1323
rect 5157 -1350 5184 -1323
rect 5220 -1350 5247 -1323
rect 2925 -1512 2961 -1476
rect 2925 -1593 2961 -1557
rect 2925 -1674 2961 -1638
rect 2925 -1755 2961 -1719
rect 2925 -2448 2961 -2412
rect 2925 -2520 2961 -2484
rect 2925 -2619 2961 -2583
rect 2925 -2691 2961 -2655
rect 3528 -2673 3555 -2646
rect 3600 -2664 3627 -2637
rect 2925 -2808 2961 -2772
rect 2925 -2889 2961 -2853
rect 2925 -2970 2961 -2934
rect 2925 -3051 2961 -3015
rect 2925 -3987 2961 -3951
rect 2925 -4059 2961 -4023
rect 2925 -4158 2961 -4122
rect 3807 -2673 3834 -2646
rect 3879 -2664 3906 -2637
rect 4212 -2646 4239 -2619
rect 4833 -2646 4860 -2619
rect 5004 -2646 5031 -2619
rect 5067 -2646 5094 -2619
rect 2925 -4230 2961 -4194
rect 3528 -4212 3555 -4185
rect 3600 -4203 3627 -4176
rect 2925 -4347 2961 -4311
rect 2925 -4428 2961 -4392
rect 2925 -4509 2961 -4473
rect 2925 -4590 2961 -4554
rect 2925 -4932 2961 -4896
rect 2925 -5004 2961 -4968
rect 2925 -5103 2961 -5067
rect 2925 -5175 2961 -5139
rect 3528 -5157 3555 -5130
rect 3600 -5148 3627 -5121
rect 2925 -5292 2961 -5256
rect 2925 -5373 2961 -5337
rect 2925 -5454 2961 -5418
rect 6633 -5220 6660 -5193
rect 6705 -5211 6732 -5184
rect 6183 -5265 6201 -5247
rect 6399 -5256 6417 -5238
rect 4833 -5301 4860 -5274
rect 5454 -5301 5481 -5274
rect 5625 -5301 5652 -5274
rect 5688 -5301 5715 -5274
rect 2925 -5535 2961 -5499
rect 2925 -5949 2961 -5913
rect 2925 -6021 2961 -5985
rect 2925 -6120 2961 -6084
rect 2925 -6192 2961 -6156
rect 3528 -6174 3555 -6147
rect 3600 -6165 3627 -6138
rect 2925 -6309 2961 -6273
rect 2925 -6390 2961 -6354
rect 2925 -6471 2961 -6435
rect 2925 -6552 2961 -6516
rect 2925 -7245 2961 -7209
rect 2925 -7317 2961 -7281
rect 2925 -7416 2961 -7380
rect 2925 -7488 2961 -7452
rect 3528 -7470 3555 -7443
rect 3600 -7461 3627 -7434
rect 2925 -7605 2961 -7569
rect 2925 -7686 2961 -7650
rect 2925 -7767 2961 -7731
rect 2925 -7848 2961 -7812
<< pdcontact >>
rect 3177 5139 3213 5175
rect 3177 5067 3213 5103
rect 3177 4968 3213 5004
rect 3528 5049 3555 5076
rect 3600 5040 3627 5067
rect 3177 4896 3213 4932
rect 3177 4779 3213 4815
rect 3177 4698 3213 4734
rect 3177 4617 3213 4653
rect 3177 4536 3213 4572
rect 4734 4779 4761 4806
rect 3897 4743 3924 4770
rect 3969 4734 3996 4761
rect 4284 4743 4302 4761
rect 4338 4734 4356 4752
rect 4437 4743 4455 4761
rect 4500 4743 4518 4761
rect 4806 4770 4833 4797
rect 3177 4194 3213 4230
rect 3177 4122 3213 4158
rect 3177 4023 3213 4059
rect 3528 4104 3555 4131
rect 3600 4095 3627 4122
rect 3177 3951 3213 3987
rect 4662 3969 4689 3996
rect 3177 3834 3213 3870
rect 3177 3753 3213 3789
rect 3879 3933 3906 3960
rect 3951 3924 3978 3951
rect 4212 3933 4230 3951
rect 4266 3924 4284 3942
rect 4365 3933 4383 3951
rect 4428 3933 4446 3951
rect 4734 3960 4761 3987
rect 5040 3933 5058 3951
rect 5094 3924 5112 3942
rect 5490 3969 5517 3996
rect 5193 3933 5211 3951
rect 5256 3933 5274 3951
rect 5562 3960 5589 3987
rect 5913 3924 5931 3942
rect 6246 3915 6264 3933
rect 6318 3924 6336 3942
rect 6372 3915 6390 3933
rect 3177 3672 3213 3708
rect 3177 3591 3213 3627
rect 3177 3177 3213 3213
rect 3177 3105 3213 3141
rect 3177 3006 3213 3042
rect 4365 3150 4392 3177
rect 4428 3141 4455 3168
rect 4491 3150 4518 3177
rect 4554 3141 4581 3168
rect 4635 3150 4662 3177
rect 4698 3141 4725 3168
rect 4761 3150 4788 3177
rect 4824 3141 4851 3168
rect 4887 3150 4914 3177
rect 4959 3141 4986 3168
rect 5157 3159 5184 3186
rect 5220 3141 5247 3168
rect 3528 3087 3555 3114
rect 3600 3078 3627 3105
rect 3861 3087 3888 3114
rect 3933 3078 3960 3105
rect 3177 2934 3213 2970
rect 3177 2817 3213 2853
rect 3177 2736 3213 2772
rect 3177 2655 3213 2691
rect 3177 2574 3213 2610
rect 3177 1881 3213 1917
rect 3177 1809 3213 1845
rect 3177 1710 3213 1746
rect 4212 1854 4239 1881
rect 4275 1845 4302 1872
rect 4338 1854 4365 1881
rect 4401 1845 4428 1872
rect 4482 1854 4509 1881
rect 4545 1845 4572 1872
rect 4608 1854 4635 1881
rect 4671 1845 4698 1872
rect 4734 1854 4761 1881
rect 4806 1845 4833 1872
rect 5004 1863 5031 1890
rect 5067 1845 5094 1872
rect 3528 1791 3555 1818
rect 3600 1782 3627 1809
rect 3807 1791 3834 1818
rect 3879 1782 3906 1809
rect 3177 1638 3213 1674
rect 3177 1521 3213 1557
rect 3177 1440 3213 1476
rect 3177 1359 3213 1395
rect 3177 1278 3213 1314
rect 3177 810 3213 846
rect 3177 738 3213 774
rect 3177 639 3213 675
rect 3528 720 3555 747
rect 3600 711 3627 738
rect 3177 567 3213 603
rect 3177 450 3213 486
rect 3177 369 3213 405
rect 3177 288 3213 324
rect 3177 207 3213 243
rect 4734 450 4761 477
rect 3897 414 3924 441
rect 3969 405 3996 432
rect 4284 414 4302 432
rect 4338 405 4356 423
rect 4437 414 4455 432
rect 4500 414 4518 432
rect 4806 441 4833 468
rect 3177 -135 3213 -99
rect 3177 -207 3213 -171
rect 3177 -306 3213 -270
rect 3528 -225 3555 -198
rect 3600 -234 3627 -207
rect 3177 -378 3213 -342
rect 4662 -360 4689 -333
rect 3177 -495 3213 -459
rect 3177 -576 3213 -540
rect 3879 -396 3906 -369
rect 3951 -405 3978 -378
rect 4212 -396 4230 -378
rect 4266 -405 4284 -387
rect 4365 -396 4383 -378
rect 4428 -396 4446 -378
rect 4734 -369 4761 -342
rect 5040 -396 5058 -378
rect 5094 -405 5112 -387
rect 5490 -360 5517 -333
rect 5193 -396 5211 -378
rect 5256 -396 5274 -378
rect 5562 -369 5589 -342
rect 5913 -405 5931 -387
rect 6246 -414 6264 -396
rect 6318 -405 6336 -387
rect 6372 -414 6390 -396
rect 3177 -657 3213 -621
rect 3177 -738 3213 -702
rect 3177 -1152 3213 -1116
rect 3177 -1224 3213 -1188
rect 3177 -1323 3213 -1287
rect 4365 -1179 4392 -1152
rect 4428 -1188 4455 -1161
rect 4491 -1179 4518 -1152
rect 4554 -1188 4581 -1161
rect 4635 -1179 4662 -1152
rect 4698 -1188 4725 -1161
rect 4761 -1179 4788 -1152
rect 4824 -1188 4851 -1161
rect 4887 -1179 4914 -1152
rect 4959 -1188 4986 -1161
rect 5157 -1170 5184 -1143
rect 5220 -1188 5247 -1161
rect 3528 -1242 3555 -1215
rect 3600 -1251 3627 -1224
rect 3861 -1242 3888 -1215
rect 3933 -1251 3960 -1224
rect 3177 -1395 3213 -1359
rect 3177 -1512 3213 -1476
rect 3177 -1593 3213 -1557
rect 3177 -1674 3213 -1638
rect 3177 -1755 3213 -1719
rect 3177 -2448 3213 -2412
rect 3177 -2520 3213 -2484
rect 3177 -2619 3213 -2583
rect 3528 -2538 3555 -2511
rect 3600 -2547 3627 -2520
rect 3177 -2691 3213 -2655
rect 3177 -2808 3213 -2772
rect 3177 -2889 3213 -2853
rect 3177 -2970 3213 -2934
rect 3177 -3051 3213 -3015
rect 3177 -3987 3213 -3951
rect 3177 -4059 3213 -4023
rect 3177 -4158 3213 -4122
rect 4212 -2475 4239 -2448
rect 4275 -2484 4302 -2457
rect 4338 -2475 4365 -2448
rect 4401 -2484 4428 -2457
rect 4482 -2475 4509 -2448
rect 4545 -2484 4572 -2457
rect 4608 -2475 4635 -2448
rect 4671 -2484 4698 -2457
rect 4734 -2475 4761 -2448
rect 4806 -2484 4833 -2457
rect 5004 -2466 5031 -2439
rect 5067 -2484 5094 -2457
rect 3807 -2538 3834 -2511
rect 3879 -2547 3906 -2520
rect 3528 -4077 3555 -4050
rect 3600 -4086 3627 -4059
rect 3177 -4230 3213 -4194
rect 3177 -4347 3213 -4311
rect 3177 -4428 3213 -4392
rect 3177 -4509 3213 -4473
rect 3177 -4590 3213 -4554
rect 3177 -4932 3213 -4896
rect 3177 -5004 3213 -4968
rect 3177 -5103 3213 -5067
rect 3528 -5022 3555 -4995
rect 3600 -5031 3627 -5004
rect 3177 -5175 3213 -5139
rect 3177 -5292 3213 -5256
rect 3177 -5373 3213 -5337
rect 3177 -5454 3213 -5418
rect 6633 -5085 6660 -5058
rect 4833 -5130 4860 -5103
rect 4896 -5139 4923 -5112
rect 4959 -5130 4986 -5103
rect 5022 -5139 5049 -5112
rect 5103 -5130 5130 -5103
rect 5166 -5139 5193 -5112
rect 5229 -5130 5256 -5103
rect 5292 -5139 5319 -5112
rect 5355 -5130 5382 -5103
rect 5427 -5139 5454 -5112
rect 5625 -5121 5652 -5094
rect 5688 -5139 5715 -5112
rect 6183 -5121 6201 -5103
rect 6237 -5130 6255 -5112
rect 6336 -5121 6354 -5103
rect 6399 -5121 6417 -5103
rect 6705 -5094 6732 -5067
rect 3177 -5535 3213 -5499
rect 3177 -5949 3213 -5913
rect 3177 -6021 3213 -5985
rect 3177 -6120 3213 -6084
rect 3528 -6039 3555 -6012
rect 3600 -6048 3627 -6021
rect 3177 -6192 3213 -6156
rect 3177 -6309 3213 -6273
rect 3177 -6390 3213 -6354
rect 3177 -6471 3213 -6435
rect 3177 -6552 3213 -6516
rect 3177 -7245 3213 -7209
rect 3177 -7317 3213 -7281
rect 3177 -7416 3213 -7380
rect 3528 -7335 3555 -7308
rect 3600 -7344 3627 -7317
rect 3177 -7488 3213 -7452
rect 3177 -7605 3213 -7569
rect 3177 -7686 3213 -7650
rect 3177 -7767 3213 -7731
rect 3177 -7848 3213 -7812
<< psubstratepcontact >>
rect 2799 4743 2835 4779
rect 2799 4653 2835 4689
rect 2799 3798 2835 3834
rect 2799 3708 2835 3744
rect 2799 2781 2835 2817
rect 2799 2691 2835 2727
rect 2799 1485 2835 1521
rect 2799 1395 2835 1431
rect 2799 414 2835 450
rect 2799 324 2835 360
rect 2799 -531 2835 -495
rect 2799 -621 2835 -585
rect 2799 -1548 2835 -1512
rect 2799 -1638 2835 -1602
rect 2799 -2844 2835 -2808
rect 2799 -2934 2835 -2898
rect 2799 -4383 2835 -4347
rect 2799 -4473 2835 -4437
rect 2799 -5328 2835 -5292
rect 2799 -5418 2835 -5382
rect 2799 -6345 2835 -6309
rect 2799 -6435 2835 -6399
rect 2799 -7641 2835 -7605
rect 2799 -7731 2835 -7695
<< nsubstratencontact >>
rect 3294 4743 3330 4779
rect 3294 4653 3330 4689
rect 3294 3798 3330 3834
rect 3294 3708 3330 3744
rect 3294 2781 3330 2817
rect 3294 2691 3330 2727
rect 3294 1485 3330 1521
rect 3294 1395 3330 1431
rect 3294 414 3330 450
rect 3294 324 3330 360
rect 3294 -531 3330 -495
rect 3294 -621 3330 -585
rect 3294 -1548 3330 -1512
rect 3294 -1638 3330 -1602
rect 3294 -2844 3330 -2808
rect 3294 -2934 3330 -2898
rect 3294 -4383 3330 -4347
rect 3294 -4473 3330 -4437
rect 3294 -5328 3330 -5292
rect 3294 -5418 3330 -5382
rect 3294 -6345 3330 -6309
rect 3294 -6435 3330 -6399
rect 3294 -7641 3330 -7605
rect 3294 -7731 3330 -7695
<< polysilicon >>
rect 2862 5220 3303 5238
rect 2862 5130 2880 5220
rect 2709 5112 2916 5130
rect 2970 5112 2979 5130
rect 2997 5112 3168 5130
rect 3231 5112 3258 5130
rect 2340 4581 2673 4599
rect 2709 4473 2727 5112
rect 2997 4959 3015 5112
rect 3285 4959 3303 5220
rect 3564 5076 3582 5094
rect 3564 4986 3582 5022
rect 2754 4941 2916 4959
rect 2970 4941 3015 4959
rect 3132 4941 3168 4959
rect 3231 4941 3303 4959
rect 3348 4959 3528 4986
rect 3573 4959 3582 4986
rect 3564 4950 3582 4959
rect 2754 4599 2772 4941
rect 3564 4905 3582 4923
rect 3042 4761 3078 4788
rect 2862 4743 2871 4761
rect 2898 4743 2916 4761
rect 2970 4743 3168 4761
rect 3231 4743 3276 4761
rect 3051 4671 3069 4743
rect 3042 4599 3078 4644
rect 2790 4581 2916 4599
rect 2970 4581 3168 4599
rect 3231 4581 3276 4599
rect 2709 4455 3078 4473
rect 3258 4392 3276 4581
rect 3600 4581 3618 4869
rect 4770 4806 4788 4923
rect 3933 4770 3951 4788
rect 4311 4770 4329 4797
rect 4473 4770 4491 4797
rect 3933 4680 3951 4716
rect 4311 4689 4329 4725
rect 3942 4653 3951 4680
rect 4023 4662 4329 4689
rect 3933 4644 3951 4653
rect 4311 4626 4329 4662
rect 4473 4653 4491 4725
rect 4770 4716 4788 4752
rect 4779 4689 4788 4716
rect 4770 4680 4788 4689
rect 4419 4635 4491 4653
rect 4770 4635 4788 4653
rect 4419 4626 4428 4635
rect 4473 4626 4491 4635
rect 3933 4599 3951 4617
rect 4311 4590 4329 4599
rect 3600 4563 3888 4581
rect 4419 4392 4428 4599
rect 4473 4590 4491 4599
rect 3258 4374 4428 4392
rect 2862 4275 3303 4293
rect 2862 4185 2880 4275
rect 2709 4167 2916 4185
rect 2970 4167 2979 4185
rect 2997 4167 3168 4185
rect 3231 4167 3258 4185
rect 2160 3636 2673 3654
rect 1872 936 2016 954
rect 1755 -4707 1773 -2043
rect 1872 -3222 1890 936
rect 2079 -693 2097 3626
rect 2709 3528 2727 4167
rect 2997 4014 3015 4167
rect 3285 4014 3303 4275
rect 3564 4131 3582 4149
rect 3564 4041 3582 4077
rect 2754 3996 2916 4014
rect 2970 3996 3015 4014
rect 3132 3996 3168 4014
rect 3231 3996 3303 4014
rect 3348 4014 3528 4041
rect 3573 4014 3582 4041
rect 3564 4005 3582 4014
rect 2754 3654 2772 3996
rect 4698 3996 4716 4113
rect 3564 3960 3582 3978
rect 3915 3960 3933 3978
rect 4239 3960 4257 3987
rect 4401 3960 4419 3987
rect 3042 3816 3078 3843
rect 2907 3798 2916 3816
rect 2970 3798 3168 3816
rect 3231 3798 3276 3816
rect 3051 3726 3069 3798
rect 3564 3771 3582 3924
rect 5067 3960 5085 3987
rect 3915 3870 3933 3906
rect 4239 3879 4257 3915
rect 3924 3843 3933 3870
rect 4023 3852 4257 3879
rect 3915 3834 3933 3843
rect 4239 3816 4257 3852
rect 4401 3843 4419 3915
rect 4698 3906 4716 3942
rect 4707 3879 4716 3906
rect 4797 3888 4914 3915
rect 4698 3870 4716 3879
rect 4887 3879 4914 3888
rect 5067 3879 5085 3915
rect 4347 3825 4419 3843
rect 4887 3852 5085 3879
rect 4698 3825 4716 3843
rect 4347 3816 4356 3825
rect 4401 3816 4419 3825
rect 5067 3816 5085 3852
rect 5157 3843 5175 4104
rect 5526 3996 5544 4113
rect 5229 3960 5247 3987
rect 5949 3951 5967 3969
rect 6003 3951 6021 4698
rect 6039 3951 6057 3969
rect 6129 3951 6147 3969
rect 6219 3951 6237 3969
rect 6345 3951 6363 3969
rect 5229 3843 5247 3915
rect 5526 3906 5544 3942
rect 5535 3879 5544 3906
rect 5526 3870 5544 3879
rect 5949 3879 5967 3906
rect 5157 3825 5247 3843
rect 6003 3879 6021 3906
rect 6039 3879 6057 3906
rect 6129 3888 6147 3906
rect 6003 3861 6057 3879
rect 5526 3825 5544 3843
rect 5229 3816 5247 3825
rect 5949 3816 5967 3861
rect 6039 3816 6057 3861
rect 6129 3816 6147 3870
rect 6219 3888 6237 3906
rect 6219 3816 6237 3870
rect 6345 3861 6363 3906
rect 6354 3843 6363 3861
rect 6345 3816 6363 3843
rect 3915 3789 3933 3807
rect 4239 3780 4257 3789
rect 3564 3753 3870 3771
rect 3042 3654 3078 3699
rect 4347 3654 4356 3789
rect 4401 3780 4419 3789
rect 5067 3780 5085 3789
rect 5229 3780 5247 3789
rect 5949 3780 5967 3789
rect 6039 3780 6057 3789
rect 6129 3780 6147 3789
rect 6219 3780 6237 3789
rect 6345 3780 6363 3789
rect 2790 3636 2916 3654
rect 2970 3636 3168 3654
rect 3231 3636 4356 3654
rect 2709 3510 3078 3528
rect 2862 3258 3303 3276
rect 2862 3168 2880 3258
rect 2709 3150 2916 3168
rect 2970 3150 2979 3168
rect 2997 3150 3168 3168
rect 3231 3150 3258 3168
rect 2151 2619 2673 2637
rect 2709 2511 2727 3150
rect 2997 2997 3015 3150
rect 3285 2997 3303 3258
rect 4401 3186 4419 3195
rect 4527 3186 4545 3195
rect 4671 3186 4689 3195
rect 4797 3186 4815 3195
rect 4932 3186 4950 3195
rect 5193 3186 5211 3195
rect 3564 3114 3582 3132
rect 3897 3114 3915 3132
rect 4401 3078 4419 3132
rect 3564 3024 3582 3060
rect 3897 3024 3915 3060
rect 4410 3051 4419 3078
rect 4527 3060 4545 3132
rect 4671 3060 4689 3132
rect 4797 3060 4815 3132
rect 4932 3060 4950 3132
rect 5193 3096 5211 3132
rect 2754 2979 2916 2997
rect 2970 2979 3015 2997
rect 3132 2979 3168 2997
rect 3231 2979 3303 2997
rect 3348 2997 3528 3024
rect 3573 2997 3582 3024
rect 3906 2997 3915 3024
rect 4401 3006 4419 3051
rect 4527 3006 4545 3033
rect 4671 3006 4689 3033
rect 4797 3006 4815 3033
rect 4932 3006 4950 3033
rect 5193 3006 5211 3069
rect 3564 2988 3582 2997
rect 3897 2988 3915 2997
rect 2754 2637 2772 2979
rect 3564 2943 3582 2961
rect 4401 2970 4419 2979
rect 4527 2970 4545 2979
rect 4671 2970 4689 2979
rect 4797 2970 4815 2979
rect 4932 2970 4950 2979
rect 5193 2970 5211 2979
rect 3897 2943 3915 2961
rect 3618 2907 3861 2925
rect 3897 2907 3906 2925
rect 3042 2799 3078 2826
rect 2853 2781 2916 2799
rect 2970 2781 3168 2799
rect 3231 2781 3276 2799
rect 3096 2718 3114 2781
rect 3042 2673 3078 2682
rect 3042 2646 3051 2673
rect 3069 2646 3078 2673
rect 3042 2637 3078 2646
rect 2790 2619 2916 2637
rect 2970 2619 3168 2637
rect 3231 2619 3276 2637
rect 2709 2493 3078 2511
rect 3123 2358 3141 2484
rect 2304 2340 3141 2358
rect 2862 1962 3303 1980
rect 2862 1872 2880 1962
rect 2709 1854 2916 1872
rect 2970 1854 2979 1872
rect 2997 1854 3168 1872
rect 3231 1854 3258 1872
rect 2709 1215 2727 1854
rect 2997 1701 3015 1854
rect 3285 1701 3303 1962
rect 4248 1890 4266 1899
rect 4374 1890 4392 1899
rect 4518 1890 4536 1899
rect 4644 1890 4662 1899
rect 4779 1890 4797 1899
rect 5040 1890 5058 1899
rect 3564 1818 3582 1836
rect 3843 1818 3861 1836
rect 4248 1782 4266 1836
rect 3564 1728 3582 1764
rect 3843 1728 3861 1764
rect 4257 1755 4266 1782
rect 4374 1764 4392 1836
rect 4518 1764 4536 1836
rect 4644 1764 4662 1836
rect 4779 1764 4797 1836
rect 5040 1800 5058 1836
rect 2754 1683 2916 1701
rect 2970 1683 3015 1701
rect 3132 1683 3168 1701
rect 3231 1683 3303 1701
rect 3348 1701 3528 1728
rect 3573 1701 3582 1728
rect 3852 1701 3861 1728
rect 4248 1710 4266 1755
rect 4374 1710 4392 1737
rect 4518 1710 4536 1737
rect 4644 1710 4662 1737
rect 4779 1710 4797 1737
rect 5040 1710 5058 1773
rect 3564 1692 3582 1701
rect 3843 1692 3861 1701
rect 2754 1341 2772 1683
rect 3564 1647 3582 1665
rect 4248 1674 4266 1683
rect 4374 1674 4392 1683
rect 4518 1674 4536 1683
rect 4644 1674 4662 1683
rect 4779 1674 4797 1683
rect 5040 1674 5058 1683
rect 3843 1647 3861 1665
rect 3042 1503 3078 1530
rect 2853 1485 2916 1503
rect 2970 1485 3168 1503
rect 3231 1485 3276 1503
rect 3096 1431 3114 1485
rect 3042 1377 3078 1386
rect 3042 1359 3051 1377
rect 3069 1359 3078 1377
rect 3042 1341 3078 1359
rect 2754 1323 2916 1341
rect 2970 1323 3168 1341
rect 3231 1323 3276 1341
rect 2709 1197 3078 1215
rect 2862 891 3303 909
rect 2862 801 2880 891
rect 2709 783 2916 801
rect 2970 783 2979 801
rect 2997 783 3168 801
rect 3231 783 3258 801
rect 2709 144 2727 783
rect 2997 630 3015 783
rect 3285 630 3303 891
rect 3429 819 3456 1440
rect 3564 747 3582 765
rect 3564 657 3582 693
rect 2754 612 2916 630
rect 2970 612 3015 630
rect 3132 612 3168 630
rect 3231 612 3303 630
rect 3348 630 3528 657
rect 3573 630 3582 657
rect 3564 621 3582 630
rect 2754 270 2772 612
rect 3564 576 3582 594
rect 3042 432 3078 459
rect 2853 414 2916 432
rect 2970 414 3168 432
rect 3231 414 3276 432
rect 3051 342 3069 414
rect 3042 270 3078 315
rect 2754 252 2916 270
rect 2970 252 3168 270
rect 3231 252 3276 270
rect 2709 126 3078 144
rect 3258 63 3276 252
rect 3600 252 3618 540
rect 4770 477 4788 594
rect 3933 441 3951 459
rect 4311 441 4329 468
rect 4473 441 4491 468
rect 3933 351 3951 387
rect 4311 360 4329 396
rect 3942 324 3951 351
rect 4023 333 4329 360
rect 3933 315 3951 324
rect 4311 297 4329 333
rect 4473 324 4491 396
rect 4770 387 4788 423
rect 4779 360 4788 387
rect 4770 351 4788 360
rect 4419 306 4491 324
rect 4770 306 4788 324
rect 4419 297 4428 306
rect 4473 297 4491 306
rect 3933 270 3951 288
rect 4311 261 4329 270
rect 3600 234 3888 252
rect 4419 63 4428 270
rect 4473 261 4491 270
rect 3258 45 4428 63
rect 3258 18 3276 45
rect 2259 0 3276 18
rect 2862 -54 3303 -36
rect 2862 -144 2880 -54
rect 2709 -162 2916 -144
rect 2970 -162 2979 -144
rect 2997 -162 3168 -144
rect 3231 -162 3258 -144
rect 2709 -801 2727 -162
rect 2997 -315 3015 -162
rect 3285 -315 3303 -54
rect 3564 -198 3582 -180
rect 3564 -288 3582 -252
rect 2754 -333 2916 -315
rect 2970 -333 3015 -315
rect 3132 -333 3168 -315
rect 3231 -333 3303 -315
rect 3348 -315 3528 -288
rect 3573 -315 3582 -288
rect 3564 -324 3582 -315
rect 2754 -675 2772 -333
rect 4698 -333 4716 -216
rect 3564 -369 3582 -351
rect 3915 -369 3933 -351
rect 4239 -369 4257 -342
rect 4401 -369 4419 -342
rect 3042 -513 3078 -486
rect 2853 -531 2916 -513
rect 2970 -531 3168 -513
rect 3231 -531 3276 -513
rect 3051 -603 3069 -531
rect 3564 -558 3582 -405
rect 5067 -369 5085 -342
rect 3915 -459 3933 -423
rect 4239 -450 4257 -414
rect 3924 -486 3933 -459
rect 4023 -477 4257 -450
rect 3915 -495 3933 -486
rect 4239 -513 4257 -477
rect 4401 -486 4419 -414
rect 4698 -423 4716 -387
rect 4707 -450 4716 -423
rect 4797 -441 4914 -414
rect 4698 -459 4716 -450
rect 4887 -450 4914 -441
rect 5067 -450 5085 -414
rect 4347 -504 4419 -486
rect 4887 -477 5085 -450
rect 4698 -504 4716 -486
rect 4347 -513 4356 -504
rect 4401 -513 4419 -504
rect 5067 -513 5085 -477
rect 5157 -486 5175 -225
rect 5526 -333 5544 -216
rect 5229 -369 5247 -342
rect 5949 -378 5967 -360
rect 6003 -378 6021 369
rect 6039 -378 6057 -360
rect 6129 -378 6147 -360
rect 6219 -378 6237 -360
rect 6345 -378 6363 -360
rect 5229 -486 5247 -414
rect 5526 -423 5544 -387
rect 5535 -450 5544 -423
rect 5526 -459 5544 -450
rect 5949 -450 5967 -423
rect 5157 -504 5247 -486
rect 6003 -450 6021 -423
rect 6039 -450 6057 -423
rect 6129 -441 6147 -423
rect 6003 -468 6057 -450
rect 5526 -504 5544 -486
rect 5229 -513 5247 -504
rect 5949 -513 5967 -468
rect 6039 -513 6057 -468
rect 6129 -513 6147 -459
rect 6219 -441 6237 -423
rect 6219 -513 6237 -459
rect 6345 -468 6363 -423
rect 6354 -486 6363 -468
rect 6345 -513 6363 -486
rect 3915 -540 3933 -522
rect 4239 -549 4257 -540
rect 3564 -576 3870 -558
rect 3042 -675 3078 -630
rect 4347 -675 4356 -540
rect 4401 -549 4419 -540
rect 5067 -549 5085 -540
rect 5229 -549 5247 -540
rect 5949 -549 5967 -540
rect 6039 -549 6057 -540
rect 6129 -549 6147 -540
rect 6219 -549 6237 -540
rect 6345 -549 6363 -540
rect 2754 -693 2799 -675
rect 2826 -693 2916 -675
rect 2970 -693 3168 -675
rect 3231 -693 4356 -675
rect 2709 -819 3078 -801
rect 2799 -990 2826 -846
rect 1953 -1008 2826 -990
rect 2862 -1071 3303 -1053
rect 2862 -1161 2880 -1071
rect 2709 -1179 2916 -1161
rect 2970 -1179 2979 -1161
rect 2997 -1179 3168 -1161
rect 3231 -1179 3258 -1161
rect 2709 -1818 2727 -1179
rect 2997 -1332 3015 -1179
rect 3285 -1332 3303 -1071
rect 4401 -1143 4419 -1134
rect 4527 -1143 4545 -1134
rect 4671 -1143 4689 -1134
rect 4797 -1143 4815 -1134
rect 4932 -1143 4950 -1134
rect 5193 -1143 5211 -1134
rect 3564 -1215 3582 -1197
rect 3897 -1215 3915 -1197
rect 4401 -1251 4419 -1197
rect 3564 -1305 3582 -1269
rect 3897 -1305 3915 -1269
rect 4410 -1278 4419 -1251
rect 4527 -1269 4545 -1197
rect 4671 -1269 4689 -1197
rect 4797 -1269 4815 -1197
rect 4932 -1269 4950 -1197
rect 5193 -1233 5211 -1197
rect 2754 -1350 2916 -1332
rect 2970 -1350 3015 -1332
rect 3132 -1350 3168 -1332
rect 3231 -1350 3303 -1332
rect 3348 -1332 3528 -1305
rect 3573 -1332 3582 -1305
rect 3906 -1332 3915 -1305
rect 4401 -1323 4419 -1278
rect 4527 -1323 4545 -1296
rect 4671 -1323 4689 -1296
rect 4797 -1323 4815 -1296
rect 4932 -1323 4950 -1296
rect 5193 -1323 5211 -1260
rect 3564 -1341 3582 -1332
rect 3897 -1341 3915 -1332
rect 2754 -1692 2772 -1350
rect 3564 -1386 3582 -1368
rect 4401 -1359 4419 -1350
rect 4527 -1359 4545 -1350
rect 4671 -1359 4689 -1350
rect 4797 -1359 4815 -1350
rect 4932 -1359 4950 -1350
rect 5193 -1359 5211 -1350
rect 3897 -1386 3915 -1368
rect 3618 -1422 3861 -1404
rect 3897 -1422 3906 -1404
rect 3042 -1530 3078 -1503
rect 2853 -1548 2916 -1530
rect 2970 -1548 3168 -1530
rect 3231 -1548 3276 -1530
rect 3096 -1611 3114 -1548
rect 3042 -1656 3078 -1647
rect 3042 -1683 3051 -1656
rect 3069 -1683 3078 -1656
rect 3042 -1692 3078 -1683
rect 2754 -1710 2799 -1692
rect 2817 -1710 2916 -1692
rect 2970 -1710 3168 -1692
rect 3231 -1710 3276 -1692
rect 2709 -1836 3078 -1818
rect 1962 -1971 1989 -1962
rect 3096 -1971 3114 -1854
rect 1962 -1989 3114 -1971
rect 1962 -6723 1989 -1989
rect 2160 -6489 2178 -2385
rect 2862 -2367 3303 -2349
rect 2862 -2457 2880 -2367
rect 2709 -2475 2916 -2457
rect 2970 -2475 2979 -2457
rect 2997 -2475 3168 -2457
rect 3231 -2475 3258 -2457
rect 2709 -3114 2727 -2475
rect 2997 -2628 3015 -2475
rect 3285 -2628 3303 -2367
rect 4248 -2439 4266 -2430
rect 4374 -2439 4392 -2430
rect 4518 -2439 4536 -2430
rect 4644 -2439 4662 -2430
rect 4779 -2439 4797 -2430
rect 5040 -2439 5058 -2430
rect 3564 -2511 3582 -2493
rect 3564 -2601 3582 -2565
rect 2754 -2646 2916 -2628
rect 2970 -2646 3015 -2628
rect 3132 -2646 3168 -2628
rect 3231 -2646 3303 -2628
rect 3348 -2628 3528 -2601
rect 3573 -2628 3582 -2601
rect 3564 -2637 3582 -2628
rect 2754 -2988 2772 -2646
rect 3564 -2682 3582 -2664
rect 3042 -2826 3078 -2799
rect 2853 -2844 2916 -2826
rect 2970 -2844 3168 -2826
rect 3231 -2844 3276 -2826
rect 3096 -2898 3114 -2844
rect 3042 -2952 3078 -2943
rect 3042 -2970 3051 -2952
rect 3069 -2970 3078 -2952
rect 3042 -2988 3078 -2970
rect 2754 -3006 2916 -2988
rect 2970 -3006 3168 -2988
rect 3231 -3006 3276 -2988
rect 2709 -3132 3078 -3114
rect 2862 -3906 3303 -3888
rect 2862 -3996 2880 -3906
rect 2709 -4014 2916 -3996
rect 2970 -4014 2979 -3996
rect 2997 -4014 3168 -3996
rect 3231 -4014 3258 -3996
rect 2709 -4653 2727 -4014
rect 2997 -4167 3015 -4014
rect 3285 -4167 3303 -3906
rect 3699 -3951 3717 -2457
rect 3843 -2511 3861 -2493
rect 4248 -2547 4266 -2493
rect 3843 -2601 3861 -2565
rect 4257 -2574 4266 -2547
rect 4374 -2565 4392 -2493
rect 4518 -2565 4536 -2493
rect 4644 -2565 4662 -2493
rect 4779 -2565 4797 -2493
rect 5040 -2529 5058 -2493
rect 3852 -2628 3861 -2601
rect 4248 -2619 4266 -2574
rect 4374 -2619 4392 -2592
rect 4518 -2619 4536 -2592
rect 4644 -2619 4662 -2592
rect 4779 -2619 4797 -2592
rect 5040 -2619 5058 -2556
rect 3843 -2637 3861 -2628
rect 4248 -2655 4266 -2646
rect 4374 -2655 4392 -2646
rect 4518 -2655 4536 -2646
rect 4644 -2655 4662 -2646
rect 4779 -2655 4797 -2646
rect 5040 -2655 5058 -2646
rect 3843 -2682 3861 -2664
rect 3564 -4050 3582 -4032
rect 3564 -4140 3582 -4104
rect 2754 -4185 2916 -4167
rect 2970 -4185 3015 -4167
rect 3132 -4185 3168 -4167
rect 3231 -4185 3303 -4167
rect 3348 -4167 3528 -4140
rect 3573 -4167 3582 -4140
rect 3654 -4158 4140 -4131
rect 3564 -4176 3582 -4167
rect 2754 -4527 2772 -4185
rect 3564 -4221 3582 -4203
rect 3042 -4365 3078 -4338
rect 2871 -4383 2916 -4365
rect 2970 -4383 3168 -4365
rect 3231 -4383 3276 -4365
rect 3042 -4527 3078 -4482
rect 2754 -4545 2916 -4527
rect 2970 -4545 3168 -4527
rect 3231 -4545 3276 -4527
rect 2709 -4671 3078 -4653
rect 3258 -4752 3276 -4545
rect 2862 -4851 3303 -4833
rect 2862 -4941 2880 -4851
rect 2709 -4959 2916 -4941
rect 2970 -4959 2979 -4941
rect 2997 -4959 3168 -4941
rect 3231 -4959 3258 -4941
rect 2709 -5598 2727 -4959
rect 2997 -5112 3015 -4959
rect 3285 -5112 3303 -4851
rect 3564 -4995 3582 -4977
rect 3564 -5085 3582 -5049
rect 2754 -5130 2916 -5112
rect 2970 -5130 3015 -5112
rect 3132 -5130 3168 -5112
rect 3231 -5130 3303 -5112
rect 3348 -5112 3528 -5085
rect 3573 -5112 3582 -5085
rect 3654 -5103 4041 -5076
rect 3564 -5121 3582 -5112
rect 2754 -5472 2772 -5130
rect 3564 -5166 3582 -5148
rect 3042 -5310 3078 -5283
rect 2871 -5328 2916 -5310
rect 2970 -5328 3168 -5310
rect 3231 -5328 3276 -5310
rect 3042 -5472 3078 -5427
rect 4023 -5427 4041 -5103
rect 4113 -5202 4140 -4158
rect 6669 -5058 6687 -4941
rect 4869 -5094 4887 -5085
rect 4995 -5094 5013 -5085
rect 5139 -5094 5157 -5085
rect 5265 -5094 5283 -5085
rect 5400 -5094 5418 -5085
rect 5661 -5094 5679 -5085
rect 6210 -5094 6228 -5067
rect 6372 -5094 6390 -5067
rect 4869 -5202 4887 -5148
rect 4113 -5229 4887 -5202
rect 4869 -5274 4887 -5229
rect 4995 -5274 5013 -5148
rect 5139 -5274 5157 -5148
rect 5265 -5274 5283 -5148
rect 5400 -5274 5418 -5148
rect 5661 -5184 5679 -5148
rect 6210 -5184 6228 -5139
rect 5769 -5211 6228 -5184
rect 5661 -5274 5679 -5211
rect 6210 -5238 6228 -5211
rect 6372 -5238 6390 -5139
rect 6669 -5148 6687 -5112
rect 6678 -5175 6687 -5148
rect 6669 -5184 6687 -5175
rect 6669 -5229 6687 -5211
rect 6210 -5274 6228 -5265
rect 6372 -5274 6390 -5265
rect 4869 -5310 4887 -5301
rect 4995 -5427 5013 -5301
rect 4023 -5454 5013 -5427
rect 2754 -5490 2916 -5472
rect 2970 -5490 3168 -5472
rect 3231 -5490 3276 -5472
rect 2709 -5616 3078 -5598
rect 3258 -5688 3276 -5490
rect 3519 -5670 4851 -5652
rect 2862 -5868 3303 -5850
rect 2862 -5958 2880 -5868
rect 2709 -5976 2916 -5958
rect 2970 -5976 2979 -5958
rect 2997 -5976 3168 -5958
rect 3231 -5976 3258 -5958
rect 2160 -6507 2673 -6489
rect 2709 -6615 2727 -5976
rect 2997 -6129 3015 -5976
rect 3285 -6129 3303 -5868
rect 3564 -6012 3582 -5994
rect 3564 -6102 3582 -6066
rect 5139 -6093 5157 -5301
rect 2754 -6147 2916 -6129
rect 2970 -6147 3015 -6129
rect 3132 -6147 3168 -6129
rect 3231 -6147 3303 -6129
rect 3348 -6129 3528 -6102
rect 3573 -6129 3582 -6102
rect 3654 -6120 5157 -6093
rect 3564 -6138 3582 -6129
rect 2754 -6489 2772 -6147
rect 3564 -6183 3582 -6165
rect 3042 -6327 3078 -6300
rect 2853 -6345 2916 -6327
rect 2970 -6345 3168 -6327
rect 3231 -6345 3276 -6327
rect 3042 -6489 3078 -6444
rect 2799 -6507 2916 -6489
rect 2970 -6507 3168 -6489
rect 3231 -6507 3249 -6489
rect 2709 -6633 3078 -6615
rect 3258 -6723 3276 -6345
rect 1962 -6741 3276 -6723
rect 2862 -7164 3303 -7146
rect 2862 -7254 2880 -7164
rect 2709 -7272 2916 -7254
rect 2970 -7272 2979 -7254
rect 2997 -7272 3168 -7254
rect 3231 -7272 3258 -7254
rect 2709 -7911 2727 -7272
rect 2997 -7425 3015 -7272
rect 3285 -7425 3303 -7164
rect 3564 -7308 3582 -7290
rect 3564 -7398 3582 -7362
rect 5265 -7389 5283 -5301
rect 5400 -5310 5418 -5301
rect 5661 -5310 5679 -5301
rect 2754 -7443 2916 -7425
rect 2970 -7443 3015 -7425
rect 3132 -7443 3168 -7425
rect 3231 -7443 3303 -7425
rect 3348 -7425 3528 -7398
rect 3573 -7425 3582 -7398
rect 3654 -7416 5283 -7389
rect 3564 -7434 3582 -7425
rect 2754 -7785 2772 -7443
rect 3564 -7479 3582 -7461
rect 3042 -7623 3078 -7596
rect 2898 -7641 2916 -7623
rect 2970 -7641 3168 -7623
rect 3231 -7641 3276 -7623
rect 3042 -7785 3078 -7740
rect 2754 -7803 2916 -7785
rect 2970 -7803 3168 -7785
rect 3231 -7803 3276 -7785
rect 2709 -7929 3078 -7911
rect 3258 -8001 3276 -7803
rect 1683 -8019 3276 -8001
<< polycontact >>
rect 2295 4581 2340 4599
rect 2673 4581 2700 4599
rect 3321 4950 3348 4986
rect 3528 4959 3573 4986
rect 3591 4869 3618 4887
rect 3042 4788 3078 4824
rect 2871 4743 2898 4761
rect 3051 4653 3069 4671
rect 2754 4581 2790 4599
rect 3042 4473 3078 4509
rect 3915 4653 3942 4680
rect 3996 4662 4023 4689
rect 4752 4689 4779 4716
rect 5994 4698 6021 4725
rect 3888 4563 3915 4581
rect 2074 3626 2099 3661
rect 2124 3636 2160 3654
rect 2673 3636 2700 3654
rect 2016 936 2052 954
rect 1755 -2043 1773 -2007
rect 3321 4005 3348 4041
rect 3528 4014 3573 4041
rect 5157 4104 5175 4158
rect 3564 3924 3582 3942
rect 3042 3843 3078 3879
rect 2871 3798 2907 3816
rect 3897 3843 3924 3870
rect 3978 3852 4023 3879
rect 4680 3879 4707 3906
rect 4761 3888 4797 3915
rect 5508 3879 5535 3906
rect 5949 3861 5967 3879
rect 6120 3870 6147 3888
rect 6219 3870 6237 3888
rect 6345 3843 6354 3861
rect 3870 3753 3915 3771
rect 3051 3708 3069 3726
rect 2754 3636 2790 3654
rect 3042 3528 3078 3564
rect 2115 2619 2151 2637
rect 2673 2619 2700 2637
rect 4383 3051 4410 3078
rect 5184 3069 5211 3096
rect 3321 2988 3348 3024
rect 3528 2997 3573 3024
rect 3879 2997 3906 3024
rect 4518 3033 4545 3060
rect 4662 3033 4689 3060
rect 4788 3033 4815 3060
rect 4923 3033 4950 3060
rect 3582 2907 3618 2925
rect 3861 2907 3897 2925
rect 3042 2826 3078 2862
rect 3096 2700 3114 2718
rect 3051 2646 3069 2673
rect 2754 2619 2790 2637
rect 3042 2511 3078 2547
rect 3123 2484 3141 2511
rect 2268 2340 2304 2358
rect 4230 1755 4257 1782
rect 5031 1773 5058 1800
rect 3321 1692 3348 1728
rect 3528 1701 3573 1728
rect 3825 1701 3852 1728
rect 4365 1737 4392 1764
rect 4509 1737 4536 1764
rect 4635 1737 4662 1764
rect 4770 1737 4797 1764
rect 3042 1530 3078 1566
rect 3429 1440 3456 1485
rect 3096 1404 3114 1431
rect 3051 1359 3069 1377
rect 3042 1215 3078 1251
rect 3429 765 3456 819
rect 3321 621 3348 657
rect 3528 630 3573 657
rect 3591 540 3618 558
rect 3042 459 3078 495
rect 3051 324 3069 342
rect 3042 144 3078 180
rect 3915 324 3942 351
rect 3996 333 4023 360
rect 4752 360 4779 387
rect 5994 369 6021 396
rect 3888 234 3915 252
rect 2187 0 2259 18
rect 2079 -729 2097 -693
rect 3321 -324 3348 -288
rect 3528 -315 3573 -288
rect 5157 -225 5175 -171
rect 3564 -405 3582 -387
rect 3042 -486 3078 -450
rect 3897 -486 3924 -459
rect 3978 -477 4023 -450
rect 4680 -450 4707 -423
rect 4761 -441 4797 -414
rect 5508 -450 5535 -423
rect 5949 -468 5967 -450
rect 6120 -459 6147 -441
rect 6219 -459 6237 -441
rect 6345 -486 6354 -468
rect 3870 -576 3915 -558
rect 3051 -621 3069 -603
rect 2799 -693 2826 -675
rect 3042 -801 3078 -765
rect 2799 -846 2826 -828
rect 1908 -1008 1953 -990
rect 4383 -1278 4410 -1251
rect 5184 -1260 5211 -1233
rect 3321 -1341 3348 -1305
rect 3528 -1332 3573 -1305
rect 3879 -1332 3906 -1305
rect 4518 -1296 4545 -1269
rect 4662 -1296 4689 -1269
rect 4788 -1296 4815 -1269
rect 4923 -1296 4950 -1269
rect 3582 -1422 3618 -1404
rect 3861 -1422 3897 -1404
rect 3042 -1503 3078 -1467
rect 3096 -1629 3114 -1611
rect 3051 -1683 3069 -1656
rect 2799 -1710 2817 -1692
rect 3042 -1818 3078 -1782
rect 3096 -1854 3114 -1818
rect 1872 -3267 1890 -3222
rect 1962 -1962 1989 -1926
rect 1755 -4734 1773 -4707
rect 2160 -2385 2178 -2340
rect 3699 -2457 3717 -2385
rect 3321 -2637 3348 -2601
rect 3528 -2628 3573 -2601
rect 3042 -2799 3078 -2763
rect 3096 -2925 3114 -2898
rect 3051 -2970 3069 -2952
rect 3042 -3114 3078 -3078
rect 4230 -2574 4257 -2547
rect 5031 -2556 5058 -2529
rect 3825 -2628 3852 -2601
rect 4365 -2592 4392 -2565
rect 4509 -2592 4536 -2565
rect 4635 -2592 4662 -2565
rect 4770 -2592 4797 -2565
rect 3699 -4041 3717 -3951
rect 3321 -4176 3348 -4140
rect 3528 -4167 3573 -4140
rect 3627 -4158 3654 -4131
rect 3042 -4338 3078 -4302
rect 2853 -4383 2871 -4365
rect 3042 -4653 3078 -4617
rect 3258 -4770 3276 -4752
rect 3321 -5121 3348 -5085
rect 3528 -5112 3573 -5085
rect 3627 -5103 3654 -5076
rect 3042 -5283 3078 -5247
rect 2853 -5328 2871 -5310
rect 5652 -5211 5679 -5184
rect 5715 -5211 5769 -5184
rect 6651 -5175 6678 -5148
rect 3042 -5598 3078 -5562
rect 3483 -5670 3519 -5652
rect 4851 -5670 4869 -5634
rect 3258 -5724 3276 -5688
rect 2673 -6507 2700 -6489
rect 3321 -6138 3348 -6102
rect 3528 -6129 3573 -6102
rect 3627 -6120 3654 -6093
rect 3042 -6300 3078 -6264
rect 2754 -6507 2799 -6489
rect 3042 -6615 3078 -6579
rect 3321 -7434 3348 -7398
rect 3528 -7425 3573 -7398
rect 3627 -7416 3654 -7389
rect 3042 -7596 3078 -7560
rect 2871 -7641 2898 -7623
rect 3042 -7911 3078 -7875
rect 1665 -8019 1683 -8001
<< metal1 >>
rect 2961 5139 3177 5175
rect 3213 5139 3393 5175
rect 2961 5067 3177 5103
rect 3213 5067 3348 5103
rect 2799 4968 2925 5004
rect 2961 4968 3177 5004
rect 3312 4986 3348 5067
rect 2799 4869 2835 4968
rect 3312 4950 3321 4986
rect 3312 4932 3348 4950
rect 2961 4896 3177 4932
rect 3213 4896 3348 4932
rect 3357 4869 3393 5139
rect 2799 4833 3024 4869
rect 2799 4779 2925 4815
rect 2799 4725 2835 4743
rect 2988 4734 3024 4833
rect 3042 4833 3393 4869
rect 3429 5130 3717 5148
rect 3042 4824 3078 4833
rect 3213 4779 3330 4815
rect 2637 4707 2835 4725
rect 2214 4581 2295 4599
rect 2637 4419 2655 4707
rect 2799 4689 2835 4707
rect 2961 4698 3177 4734
rect 3294 4725 3330 4743
rect 3429 4725 3456 5130
rect 3519 5121 3555 5130
rect 3528 5076 3555 5121
rect 3600 4995 3627 5040
rect 3600 4968 3663 4995
rect 3600 4950 3627 4968
rect 3528 4887 3555 4914
rect 3294 4698 3456 4725
rect 3501 4869 3591 4887
rect 3294 4689 3330 4698
rect 3069 4653 3096 4671
rect 2799 4617 2925 4653
rect 3213 4617 3330 4653
rect 2700 4581 2754 4599
rect 2961 4536 3177 4572
rect 3042 4509 3078 4536
rect 3501 4419 3519 4869
rect 2637 4401 3519 4419
rect 3699 4833 3717 5130
rect 4734 4860 4833 4869
rect 4734 4833 4761 4860
rect 3699 4815 4761 4833
rect 2421 4329 2574 4347
rect 1674 3798 2322 3816
rect 1674 -990 1701 3798
rect 2637 3780 2655 4401
rect 2961 4194 3177 4230
rect 3213 4194 3393 4230
rect 3699 4203 3717 4815
rect 3897 4770 3924 4815
rect 4284 4761 4302 4815
rect 4437 4761 4455 4815
rect 4734 4806 4761 4815
rect 3969 4644 3996 4734
rect 4338 4680 4356 4734
rect 4500 4680 4518 4743
rect 4806 4725 4833 4770
rect 4662 4689 4752 4716
rect 4806 4698 5994 4725
rect 4662 4680 4680 4689
rect 4338 4662 4680 4680
rect 4806 4680 4833 4698
rect 4500 4626 4518 4662
rect 3897 4581 3924 4608
rect 4734 4617 4761 4644
rect 4284 4581 4302 4599
rect 4734 4599 4833 4617
rect 4734 4581 4770 4599
rect 3915 4563 4770 4581
rect 2961 4122 3177 4158
rect 3213 4122 3348 4158
rect 2799 4023 2925 4059
rect 2961 4023 3177 4059
rect 3312 4041 3348 4122
rect 2799 3924 2835 4023
rect 3312 4005 3321 4041
rect 3312 3987 3348 4005
rect 2961 3951 3177 3987
rect 3213 3951 3348 3987
rect 3357 3924 3393 4194
rect 2799 3888 3024 3924
rect 2799 3834 2925 3870
rect 2799 3780 2835 3798
rect 2988 3789 3024 3888
rect 3042 3888 3393 3924
rect 3429 4185 3717 4203
rect 3042 3879 3078 3888
rect 3213 3834 3330 3870
rect 2637 3762 2835 3780
rect 2099 3636 2124 3654
rect 2637 3474 2655 3762
rect 2799 3744 2835 3762
rect 2961 3753 3177 3789
rect 3294 3780 3330 3798
rect 3429 3780 3456 4185
rect 3519 4176 3555 4185
rect 3528 4131 3555 4176
rect 3600 4050 3627 4095
rect 3600 4023 3654 4050
rect 3699 4023 3717 4185
rect 5157 4158 5175 4248
rect 4662 4050 4761 4059
rect 5490 4050 5931 4068
rect 4662 4023 4689 4050
rect 5490 4023 5517 4050
rect 3600 4005 3627 4023
rect 3699 4005 5517 4023
rect 3528 3942 3555 3969
rect 3294 3753 3456 3780
rect 3501 3924 3564 3942
rect 3582 3924 3618 3942
rect 3294 3744 3330 3753
rect 3069 3708 3096 3726
rect 2799 3672 2925 3708
rect 3213 3672 3330 3708
rect 2700 3636 2754 3654
rect 2961 3591 3177 3627
rect 3042 3564 3078 3591
rect 3501 3474 3519 3924
rect 2637 3456 3519 3474
rect 2637 2763 2655 3456
rect 3699 3249 3717 4005
rect 3879 3960 3906 4005
rect 4212 3951 4230 4005
rect 4365 3951 4383 4005
rect 4662 3996 4689 4005
rect 3951 3834 3978 3924
rect 4266 3870 4284 3924
rect 4428 3870 4446 3933
rect 4590 3879 4680 3906
rect 4590 3870 4608 3879
rect 4266 3852 4608 3870
rect 4734 3870 4761 3960
rect 5040 3951 5058 4005
rect 5193 3951 5211 4005
rect 5490 3996 5517 4005
rect 5913 3996 5931 4050
rect 4428 3816 4446 3852
rect 3879 3771 3906 3798
rect 5094 3870 5112 3924
rect 5256 3870 5274 3933
rect 5562 3915 5589 3960
rect 5913 3978 6363 3996
rect 5913 3942 5931 3978
rect 6318 3942 6336 3978
rect 5418 3879 5508 3906
rect 5562 3888 5769 3915
rect 5418 3870 5436 3879
rect 5094 3852 5436 3870
rect 5562 3870 5589 3888
rect 4662 3807 4689 3834
rect 5256 3816 5274 3852
rect 4212 3771 4230 3789
rect 4662 3789 4761 3807
rect 5751 3879 5769 3888
rect 5751 3861 5949 3879
rect 6246 3861 6264 3915
rect 6372 3861 6390 3915
rect 5976 3843 6345 3861
rect 6372 3843 6417 3861
rect 5490 3807 5517 3834
rect 5976 3816 5994 3843
rect 6066 3816 6084 3843
rect 6156 3816 6174 3843
rect 6246 3816 6264 3843
rect 6372 3816 6390 3843
rect 4662 3771 4698 3789
rect 5040 3771 5058 3789
rect 5490 3789 5589 3807
rect 5490 3771 5526 3789
rect 5913 3771 5931 3798
rect 6012 3771 6030 3798
rect 6102 3771 6120 3798
rect 6192 3771 6210 3798
rect 6318 3771 6336 3798
rect 3915 3753 6336 3771
rect 3699 3222 5193 3249
rect 2961 3177 3177 3213
rect 3213 3177 3393 3213
rect 3699 3186 3717 3222
rect 2961 3105 3177 3141
rect 3213 3105 3348 3141
rect 2799 3006 2925 3042
rect 2961 3006 3177 3042
rect 3312 3024 3348 3105
rect 2799 2907 2835 3006
rect 3312 2988 3321 3024
rect 3312 2970 3348 2988
rect 2961 2934 3177 2970
rect 3213 2934 3348 2970
rect 3357 2907 3393 3177
rect 2799 2871 3024 2907
rect 2799 2817 2925 2853
rect 2799 2763 2835 2781
rect 2988 2772 3024 2871
rect 3042 2871 3393 2907
rect 3429 3177 3717 3186
rect 4365 3177 4392 3222
rect 3429 3168 3960 3177
rect 3042 2862 3078 2871
rect 3213 2817 3330 2853
rect 2637 2745 2835 2763
rect 1962 2619 2115 2637
rect 1674 -1008 1908 -990
rect 1755 -2007 1773 -1926
rect 1620 -2133 1728 -2106
rect 1755 -4788 1773 -4734
rect 1809 -5733 1827 -1008
rect 1962 -1926 1989 2619
rect 2637 2457 2655 2745
rect 2799 2727 2835 2745
rect 2961 2736 3177 2772
rect 3294 2763 3330 2781
rect 3429 2763 3456 3168
rect 3519 3159 3555 3168
rect 3528 3114 3555 3159
rect 3699 3159 3888 3168
rect 3600 2988 3627 3078
rect 3528 2925 3555 2952
rect 3294 2736 3456 2763
rect 3501 2907 3582 2925
rect 3294 2727 3330 2736
rect 2799 2655 2925 2691
rect 3096 2682 3114 2700
rect 3213 2655 3330 2691
rect 2700 2619 2754 2637
rect 2961 2574 3177 2610
rect 3042 2547 3078 2574
rect 3123 2511 3141 2529
rect 3501 2457 3519 2907
rect 2637 2439 3519 2457
rect 2250 2340 2268 2358
rect 2331 2277 2556 2295
rect 2637 1467 2655 2439
rect 3699 1953 3717 3159
rect 3861 3114 3888 3159
rect 4491 3177 4518 3222
rect 4635 3177 4662 3222
rect 4428 3096 4455 3141
rect 4761 3177 4788 3222
rect 4554 3096 4581 3141
rect 4887 3177 4914 3222
rect 4698 3096 4725 3141
rect 5157 3186 5184 3222
rect 4824 3096 4851 3141
rect 4959 3096 4986 3141
rect 5220 3096 5247 3141
rect 6093 3096 6111 3447
rect 3933 3033 3960 3078
rect 4158 3051 4383 3078
rect 4428 3069 5184 3096
rect 5220 3069 6111 3096
rect 4158 3033 4176 3051
rect 4761 3033 4788 3060
rect 3933 3006 4176 3033
rect 4986 3006 5013 3069
rect 5220 3006 5247 3069
rect 3933 2988 3960 3006
rect 3861 2925 3888 2952
rect 4365 2934 4392 2979
rect 5157 2934 5184 2979
rect 4365 2925 5184 2934
rect 3852 2907 3861 2925
rect 3897 2907 5184 2925
rect 3699 1926 5040 1953
rect 2961 1881 3177 1917
rect 3213 1881 3393 1917
rect 3699 1890 3717 1926
rect 2961 1809 3177 1845
rect 3213 1809 3348 1845
rect 2799 1710 2925 1746
rect 2961 1710 3177 1746
rect 3312 1728 3348 1809
rect 2799 1611 2835 1710
rect 3312 1692 3321 1728
rect 3312 1674 3348 1692
rect 2961 1638 3177 1674
rect 3213 1638 3348 1674
rect 3357 1611 3393 1881
rect 2799 1575 3024 1611
rect 2799 1521 2925 1557
rect 2799 1467 2835 1485
rect 2988 1476 3024 1575
rect 3042 1575 3393 1611
rect 3429 1872 3906 1890
rect 4212 1881 4239 1926
rect 3042 1566 3078 1575
rect 3213 1521 3330 1557
rect 2637 1449 2835 1467
rect 2637 1161 2655 1449
rect 2799 1431 2835 1449
rect 2961 1440 3177 1476
rect 3294 1467 3330 1485
rect 3429 1485 3456 1872
rect 3519 1863 3555 1872
rect 3798 1863 3834 1872
rect 3528 1818 3555 1863
rect 3807 1818 3834 1863
rect 4338 1881 4365 1926
rect 4482 1881 4509 1926
rect 3600 1737 3627 1782
rect 4275 1800 4302 1845
rect 4608 1881 4635 1926
rect 4401 1800 4428 1845
rect 4734 1881 4761 1926
rect 4545 1800 4572 1845
rect 5004 1890 5031 1926
rect 4671 1800 4698 1845
rect 4806 1800 4833 1845
rect 5067 1800 5094 1845
rect 6183 1800 6201 3033
rect 3879 1737 3906 1782
rect 4068 1755 4230 1782
rect 4275 1773 5031 1800
rect 5067 1773 6201 1800
rect 4068 1737 4086 1755
rect 3600 1710 3654 1737
rect 3600 1692 3627 1710
rect 3879 1710 4086 1737
rect 4833 1710 4860 1773
rect 5067 1710 5094 1773
rect 3879 1692 3906 1710
rect 3528 1629 3555 1656
rect 3807 1629 3834 1656
rect 4212 1638 4239 1683
rect 5004 1638 5031 1683
rect 4212 1629 5031 1638
rect 3294 1440 3429 1467
rect 3501 1611 5031 1629
rect 3294 1431 3330 1440
rect 3096 1395 3114 1404
rect 2799 1359 2925 1395
rect 3213 1359 3330 1395
rect 2961 1278 3177 1314
rect 3042 1251 3078 1278
rect 3501 1161 3519 1611
rect 2637 1143 3519 1161
rect 2250 1017 2277 1035
rect 2052 936 2241 954
rect 2637 396 2655 1143
rect 3249 1044 3267 1053
rect 2961 810 3177 846
rect 3213 810 3393 846
rect 2961 738 3177 774
rect 3213 738 3348 774
rect 2799 639 2925 675
rect 2961 639 3177 675
rect 3312 657 3348 738
rect 2799 540 2835 639
rect 3312 621 3321 657
rect 3312 603 3348 621
rect 2961 567 3177 603
rect 3213 567 3348 603
rect 3357 540 3393 810
rect 2799 504 3024 540
rect 2799 450 2925 486
rect 2799 396 2835 414
rect 2988 405 3024 504
rect 3042 504 3393 540
rect 3456 801 3717 819
rect 3519 792 3555 801
rect 3042 495 3078 504
rect 3213 450 3330 486
rect 2637 378 2835 396
rect 2637 90 2655 378
rect 2799 360 2835 378
rect 2961 369 3177 405
rect 3294 396 3330 414
rect 3429 396 3456 765
rect 3528 747 3555 792
rect 3600 666 3627 711
rect 3600 639 3663 666
rect 3600 621 3627 639
rect 3528 558 3555 585
rect 3294 369 3456 396
rect 3501 540 3591 558
rect 3294 360 3330 369
rect 3069 324 3096 342
rect 2799 288 2925 324
rect 3213 288 3330 324
rect 2961 207 3177 243
rect 3042 180 3078 207
rect 3501 90 3519 540
rect 2637 72 3519 90
rect 3699 504 3717 801
rect 4734 531 4833 540
rect 4734 504 4761 531
rect 3699 486 4761 504
rect 2160 0 2187 18
rect 2637 -549 2655 72
rect 2961 -135 3177 -99
rect 3213 -135 3393 -99
rect 3699 -126 3717 486
rect 3897 441 3924 486
rect 4284 432 4302 486
rect 4437 432 4455 486
rect 4734 477 4761 486
rect 3969 315 3996 405
rect 4338 351 4356 405
rect 4500 351 4518 414
rect 4806 396 4833 441
rect 4662 360 4752 387
rect 4806 369 5994 396
rect 4662 351 4680 360
rect 4338 333 4680 351
rect 4806 351 4833 369
rect 4500 297 4518 333
rect 3897 252 3924 279
rect 4734 288 4761 315
rect 4284 252 4302 270
rect 4734 270 4833 288
rect 4734 252 4770 270
rect 3915 234 4770 252
rect 2961 -207 3177 -171
rect 3213 -207 3348 -171
rect 2799 -306 2925 -270
rect 2961 -306 3177 -270
rect 3312 -288 3348 -207
rect 2799 -405 2835 -306
rect 3312 -324 3321 -288
rect 3312 -342 3348 -324
rect 2961 -378 3177 -342
rect 3213 -378 3348 -342
rect 3357 -405 3393 -135
rect 2799 -441 3024 -405
rect 2799 -495 2925 -459
rect 2799 -549 2835 -531
rect 2988 -540 3024 -441
rect 3042 -441 3393 -405
rect 3429 -144 3717 -126
rect 3042 -450 3078 -441
rect 3213 -495 3330 -459
rect 2637 -567 2835 -549
rect 2079 -936 2097 -729
rect 2637 -855 2655 -567
rect 2799 -585 2835 -567
rect 2961 -576 3177 -540
rect 3294 -549 3330 -531
rect 3429 -549 3456 -144
rect 3519 -153 3555 -144
rect 3528 -198 3555 -153
rect 3600 -279 3627 -234
rect 3600 -306 3654 -279
rect 3699 -306 3717 -144
rect 5157 -171 5175 -81
rect 4662 -279 4761 -270
rect 5490 -279 5931 -261
rect 4662 -306 4689 -279
rect 5490 -306 5517 -279
rect 3600 -324 3627 -306
rect 3699 -324 5517 -306
rect 3528 -387 3555 -360
rect 3294 -576 3456 -549
rect 3501 -405 3564 -387
rect 3582 -405 3618 -387
rect 3294 -585 3330 -576
rect 3069 -621 3096 -603
rect 2799 -657 2925 -621
rect 3213 -657 3330 -621
rect 2799 -828 2826 -693
rect 2961 -738 3177 -702
rect 3042 -765 3078 -738
rect 3501 -855 3519 -405
rect 1872 -3285 1890 -3267
rect 2079 -5697 2097 -954
rect 2160 -2340 2178 -2133
rect 2196 -4743 2214 -891
rect 2637 -873 3519 -855
rect 2637 -1566 2655 -873
rect 3699 -1080 3717 -324
rect 3879 -369 3906 -324
rect 4212 -378 4230 -324
rect 4365 -378 4383 -324
rect 4662 -333 4689 -324
rect 3871 -486 3879 -459
rect 3951 -495 3978 -405
rect 4266 -459 4284 -405
rect 4428 -459 4446 -396
rect 4590 -450 4680 -423
rect 4590 -459 4608 -450
rect 4266 -477 4608 -459
rect 4734 -459 4761 -369
rect 5040 -378 5058 -324
rect 5193 -378 5211 -324
rect 5490 -333 5517 -324
rect 5913 -333 5931 -279
rect 4428 -513 4446 -477
rect 3879 -558 3906 -531
rect 5094 -459 5112 -405
rect 5256 -459 5274 -396
rect 5562 -414 5589 -369
rect 5913 -351 6363 -333
rect 5913 -387 5931 -351
rect 6318 -387 6336 -351
rect 5418 -450 5508 -423
rect 5562 -441 5769 -414
rect 5418 -459 5436 -450
rect 5094 -477 5436 -459
rect 5562 -459 5589 -441
rect 4662 -522 4689 -495
rect 5256 -513 5274 -477
rect 4212 -558 4230 -540
rect 4662 -540 4761 -522
rect 5751 -450 5769 -441
rect 5751 -468 5949 -450
rect 6246 -468 6264 -414
rect 6372 -468 6390 -414
rect 5976 -486 6345 -468
rect 6372 -486 6417 -468
rect 5490 -522 5517 -495
rect 5976 -513 5994 -486
rect 6066 -513 6084 -486
rect 6156 -513 6174 -486
rect 6246 -513 6264 -486
rect 6372 -513 6390 -486
rect 4662 -558 4698 -540
rect 5040 -558 5058 -540
rect 5490 -540 5589 -522
rect 5490 -558 5526 -540
rect 5913 -558 5931 -531
rect 6012 -558 6030 -531
rect 6102 -558 6120 -531
rect 6192 -558 6210 -531
rect 6318 -558 6336 -531
rect 3915 -576 6336 -558
rect 3699 -1107 5193 -1080
rect 2961 -1152 3177 -1116
rect 3213 -1152 3393 -1116
rect 3699 -1143 3717 -1107
rect 2961 -1224 3177 -1188
rect 3213 -1224 3348 -1188
rect 2799 -1323 2925 -1287
rect 2961 -1323 3177 -1287
rect 3312 -1305 3348 -1224
rect 2799 -1422 2835 -1323
rect 3312 -1341 3321 -1305
rect 3312 -1359 3348 -1341
rect 2961 -1395 3177 -1359
rect 3213 -1395 3348 -1359
rect 3357 -1422 3393 -1152
rect 2799 -1458 3024 -1422
rect 2799 -1512 2925 -1476
rect 2799 -1566 2835 -1548
rect 2988 -1557 3024 -1458
rect 3042 -1458 3393 -1422
rect 3429 -1152 3717 -1143
rect 4365 -1152 4392 -1107
rect 3429 -1161 3960 -1152
rect 3042 -1467 3078 -1458
rect 3213 -1512 3330 -1476
rect 2637 -1584 2835 -1566
rect 2637 -1872 2655 -1584
rect 2799 -1602 2835 -1584
rect 2961 -1593 3177 -1557
rect 3294 -1566 3330 -1548
rect 3429 -1566 3456 -1161
rect 3519 -1170 3555 -1161
rect 3528 -1215 3555 -1170
rect 3699 -1170 3888 -1161
rect 3600 -1341 3627 -1251
rect 3528 -1404 3555 -1377
rect 3294 -1593 3456 -1566
rect 3501 -1422 3582 -1404
rect 3294 -1602 3330 -1593
rect 2799 -1674 2925 -1638
rect 3096 -1647 3114 -1629
rect 3213 -1674 3330 -1638
rect 2799 -1728 2817 -1710
rect 2961 -1755 3177 -1719
rect 3042 -1782 3078 -1755
rect 3096 -1818 3114 -1800
rect 3501 -1872 3519 -1422
rect 2637 -1890 3519 -1872
rect 2637 -2862 2655 -1890
rect 3699 -2376 3717 -1170
rect 3861 -1215 3888 -1170
rect 4491 -1152 4518 -1107
rect 4635 -1152 4662 -1107
rect 4428 -1233 4455 -1188
rect 4761 -1152 4788 -1107
rect 4554 -1233 4581 -1188
rect 4887 -1152 4914 -1107
rect 4698 -1233 4725 -1188
rect 5157 -1143 5184 -1107
rect 4824 -1233 4851 -1188
rect 4959 -1233 4986 -1188
rect 5220 -1233 5247 -1188
rect 6093 -1233 6111 -882
rect 3933 -1296 3960 -1251
rect 4158 -1278 4383 -1251
rect 4428 -1260 5184 -1233
rect 5220 -1260 6111 -1233
rect 4158 -1296 4176 -1278
rect 4761 -1296 4788 -1269
rect 3933 -1323 4176 -1296
rect 4986 -1323 5013 -1260
rect 5220 -1323 5247 -1260
rect 3933 -1341 3960 -1323
rect 3861 -1404 3888 -1377
rect 4365 -1395 4392 -1350
rect 5157 -1395 5184 -1350
rect 4365 -1404 5184 -1395
rect 3852 -1422 3861 -1404
rect 3897 -1422 5184 -1404
rect 3699 -2385 5040 -2376
rect 2961 -2448 3177 -2412
rect 3213 -2448 3393 -2412
rect 2961 -2520 3177 -2484
rect 3213 -2520 3348 -2484
rect 2799 -2619 2925 -2583
rect 2961 -2619 3177 -2583
rect 3312 -2601 3348 -2520
rect 2799 -2718 2835 -2619
rect 3312 -2637 3321 -2601
rect 3312 -2655 3348 -2637
rect 2961 -2691 3177 -2655
rect 3213 -2691 3348 -2655
rect 3357 -2718 3393 -2448
rect 2799 -2754 3024 -2718
rect 2799 -2808 2925 -2772
rect 2799 -2862 2835 -2844
rect 2988 -2853 3024 -2754
rect 3042 -2754 3393 -2718
rect 3429 -2457 3699 -2439
rect 3717 -2403 5040 -2385
rect 3717 -2457 3906 -2439
rect 4212 -2448 4239 -2403
rect 3042 -2763 3078 -2754
rect 3213 -2808 3330 -2772
rect 2637 -2880 2835 -2862
rect 2637 -3168 2655 -2880
rect 2799 -2898 2835 -2880
rect 2961 -2889 3177 -2853
rect 3294 -2862 3330 -2844
rect 3429 -2862 3456 -2457
rect 3519 -2466 3555 -2457
rect 3798 -2466 3834 -2457
rect 3528 -2511 3555 -2466
rect 3807 -2511 3834 -2466
rect 4338 -2448 4365 -2403
rect 4482 -2448 4509 -2403
rect 3600 -2592 3627 -2547
rect 4275 -2529 4302 -2484
rect 4608 -2448 4635 -2403
rect 4401 -2529 4428 -2484
rect 4734 -2448 4761 -2403
rect 4545 -2529 4572 -2484
rect 5004 -2439 5031 -2403
rect 4671 -2529 4698 -2484
rect 4806 -2529 4833 -2484
rect 5067 -2529 5094 -2484
rect 6183 -2529 6201 -1296
rect 3879 -2592 3906 -2547
rect 4068 -2574 4230 -2547
rect 4275 -2556 5031 -2529
rect 5067 -2556 6201 -2529
rect 4068 -2592 4086 -2574
rect 3600 -2619 3654 -2592
rect 3600 -2637 3627 -2619
rect 3879 -2619 4086 -2592
rect 4833 -2619 4860 -2556
rect 5067 -2619 5094 -2556
rect 3879 -2637 3906 -2619
rect 3528 -2700 3555 -2673
rect 3807 -2700 3834 -2673
rect 4212 -2691 4239 -2646
rect 5004 -2691 5031 -2646
rect 4212 -2700 5031 -2691
rect 3294 -2889 3456 -2862
rect 3501 -2718 5031 -2700
rect 3294 -2898 3330 -2889
rect 3096 -2934 3114 -2925
rect 2799 -2970 2925 -2934
rect 3213 -2970 3330 -2934
rect 2961 -3051 3177 -3015
rect 3042 -3078 3078 -3051
rect 3501 -3168 3519 -2718
rect 2637 -3186 3519 -3168
rect 2637 -4401 2655 -3186
rect 2961 -3987 3177 -3951
rect 3213 -3987 3393 -3951
rect 2961 -4059 3177 -4023
rect 3213 -4059 3348 -4023
rect 2799 -4158 2925 -4122
rect 2961 -4158 3177 -4122
rect 3312 -4140 3348 -4059
rect 2799 -4257 2835 -4158
rect 3312 -4176 3321 -4140
rect 3312 -4194 3348 -4176
rect 2961 -4230 3177 -4194
rect 3213 -4230 3348 -4194
rect 3357 -4257 3393 -3987
rect 2799 -4293 3024 -4257
rect 2799 -4347 2925 -4311
rect 2799 -4401 2835 -4383
rect 2637 -4419 2835 -4401
rect 2637 -4707 2655 -4419
rect 2799 -4437 2835 -4419
rect 2853 -4401 2871 -4383
rect 2988 -4392 3024 -4293
rect 3042 -4293 3393 -4257
rect 3429 -3996 3699 -3978
rect 3042 -4302 3078 -4293
rect 3213 -4347 3330 -4311
rect 2961 -4428 3177 -4392
rect 3294 -4401 3330 -4383
rect 3429 -4401 3456 -3996
rect 3519 -4005 3555 -3996
rect 3528 -4050 3555 -4005
rect 3600 -4176 3627 -4086
rect 3528 -4239 3555 -4212
rect 3294 -4428 3456 -4401
rect 3501 -4257 3618 -4239
rect 3294 -4437 3330 -4428
rect 2799 -4509 2925 -4473
rect 3213 -4509 3330 -4473
rect 2961 -4590 3177 -4554
rect 3042 -4617 3078 -4590
rect 3501 -4707 3519 -4257
rect 2637 -4725 3519 -4707
rect 2637 -5346 2655 -4725
rect 3258 -4788 3276 -4770
rect 2961 -4932 3177 -4896
rect 3213 -4932 3393 -4896
rect 3699 -4923 3717 -4041
rect 2961 -5004 3177 -4968
rect 3213 -5004 3348 -4968
rect 2799 -5103 2925 -5067
rect 2961 -5103 3177 -5067
rect 3312 -5085 3348 -5004
rect 2799 -5202 2835 -5103
rect 3312 -5121 3321 -5085
rect 3312 -5139 3348 -5121
rect 2961 -5175 3177 -5139
rect 3213 -5175 3348 -5139
rect 3357 -5202 3393 -4932
rect 2799 -5238 3024 -5202
rect 2799 -5292 2925 -5256
rect 2799 -5346 2835 -5328
rect 2637 -5364 2835 -5346
rect 2637 -5652 2655 -5364
rect 2799 -5382 2835 -5364
rect 2853 -5346 2871 -5328
rect 2988 -5337 3024 -5238
rect 3042 -5238 3393 -5202
rect 3429 -4941 4860 -4923
rect 3042 -5247 3078 -5238
rect 3213 -5292 3330 -5256
rect 2961 -5373 3177 -5337
rect 3294 -5346 3330 -5328
rect 3429 -5346 3456 -4941
rect 3519 -4950 3555 -4941
rect 3528 -4995 3555 -4950
rect 3600 -5121 3627 -5031
rect 3528 -5184 3555 -5157
rect 3294 -5373 3456 -5346
rect 3501 -5202 3618 -5184
rect 3294 -5382 3330 -5373
rect 2799 -5454 2925 -5418
rect 3213 -5454 3330 -5418
rect 2961 -5535 3177 -5499
rect 3042 -5562 3078 -5535
rect 3501 -5652 3519 -5202
rect 2637 -5670 3483 -5652
rect 2637 -6363 2655 -5670
rect 3258 -5733 3276 -5724
rect 2961 -5949 3177 -5913
rect 3213 -5949 3393 -5913
rect 3699 -5940 3717 -4941
rect 4833 -5031 4860 -4941
rect 6633 -5004 6732 -4995
rect 6633 -5031 6660 -5004
rect 4833 -5049 6660 -5031
rect 4833 -5058 5661 -5049
rect 4833 -5103 4860 -5058
rect 4959 -5103 4986 -5058
rect 5103 -5103 5130 -5058
rect 4896 -5184 4923 -5139
rect 5229 -5103 5256 -5058
rect 5022 -5184 5049 -5139
rect 5355 -5103 5382 -5058
rect 5166 -5184 5193 -5139
rect 5625 -5094 5652 -5058
rect 5292 -5184 5319 -5139
rect 6183 -5103 6201 -5049
rect 5427 -5184 5454 -5139
rect 6336 -5103 6354 -5049
rect 6633 -5058 6660 -5049
rect 4896 -5211 5652 -5184
rect 5454 -5274 5481 -5211
rect 5688 -5274 5715 -5139
rect 6237 -5184 6255 -5130
rect 6399 -5184 6417 -5121
rect 6705 -5139 6732 -5094
rect 6561 -5175 6651 -5148
rect 6705 -5166 6759 -5139
rect 6561 -5184 6579 -5175
rect 6237 -5202 6579 -5184
rect 6705 -5184 6732 -5166
rect 6399 -5238 6417 -5202
rect 6633 -5247 6660 -5220
rect 6183 -5283 6201 -5265
rect 6633 -5265 6732 -5247
rect 6633 -5283 6669 -5265
rect 6183 -5301 6669 -5283
rect 4833 -5346 4860 -5301
rect 5625 -5346 5652 -5301
rect 6201 -5346 6219 -5301
rect 4833 -5373 6219 -5346
rect 4851 -5634 4869 -5373
rect 2961 -6021 3177 -5985
rect 3213 -6021 3348 -5985
rect 2799 -6120 2925 -6084
rect 2961 -6120 3177 -6084
rect 3312 -6102 3348 -6021
rect 2799 -6219 2835 -6120
rect 3312 -6138 3321 -6102
rect 3312 -6156 3348 -6138
rect 2961 -6192 3177 -6156
rect 3213 -6192 3348 -6156
rect 3357 -6219 3393 -5949
rect 2799 -6255 3024 -6219
rect 2799 -6309 2925 -6273
rect 2799 -6363 2835 -6345
rect 2988 -6354 3024 -6255
rect 3042 -6255 3393 -6219
rect 3429 -5958 3717 -5940
rect 3042 -6264 3078 -6255
rect 3213 -6309 3330 -6273
rect 2637 -6381 2835 -6363
rect 2637 -6669 2655 -6381
rect 2799 -6399 2835 -6381
rect 2961 -6390 3177 -6354
rect 3294 -6363 3330 -6345
rect 3429 -6363 3456 -5958
rect 3519 -5967 3555 -5958
rect 3528 -6012 3555 -5967
rect 3600 -6138 3627 -6048
rect 3528 -6201 3555 -6174
rect 3294 -6390 3456 -6363
rect 3501 -6219 3618 -6201
rect 3294 -6399 3330 -6390
rect 2799 -6471 2925 -6435
rect 3213 -6471 3330 -6435
rect 2700 -6507 2754 -6489
rect 2961 -6552 3177 -6516
rect 3042 -6579 3078 -6552
rect 3501 -6669 3519 -6219
rect 2637 -6687 3519 -6669
rect 2637 -7659 2655 -6687
rect 2961 -7245 3177 -7209
rect 3213 -7245 3393 -7209
rect 3699 -7236 3717 -5958
rect 2961 -7317 3177 -7281
rect 3213 -7317 3348 -7281
rect 2799 -7416 2925 -7380
rect 2961 -7416 3177 -7380
rect 3312 -7398 3348 -7317
rect 2799 -7515 2835 -7416
rect 3312 -7434 3321 -7398
rect 3312 -7452 3348 -7434
rect 2961 -7488 3177 -7452
rect 3213 -7488 3348 -7452
rect 3357 -7515 3393 -7245
rect 2799 -7551 3024 -7515
rect 2799 -7605 2925 -7569
rect 2799 -7659 2835 -7641
rect 2988 -7650 3024 -7551
rect 3042 -7551 3393 -7515
rect 3429 -7254 3717 -7236
rect 3042 -7560 3078 -7551
rect 3213 -7605 3330 -7569
rect 2637 -7677 2835 -7659
rect 2637 -7965 2655 -7677
rect 2799 -7695 2835 -7677
rect 2961 -7686 3177 -7650
rect 3294 -7659 3330 -7641
rect 3429 -7659 3456 -7254
rect 3519 -7263 3555 -7254
rect 3528 -7308 3555 -7263
rect 3600 -7434 3627 -7344
rect 3528 -7497 3555 -7470
rect 3294 -7686 3456 -7659
rect 3501 -7515 3618 -7497
rect 3294 -7695 3330 -7686
rect 2799 -7767 2925 -7731
rect 3213 -7767 3330 -7731
rect 2961 -7848 3177 -7812
rect 3042 -7875 3078 -7848
rect 3501 -7965 3519 -7515
rect 2637 -7983 3519 -7965
rect 1665 -8001 1683 -7983
<< m2contact >>
rect 2844 4743 2871 4761
rect 2196 4572 2214 4599
rect 3096 4653 3114 4671
rect 2322 3798 2367 3816
rect 3888 4653 3915 4680
rect 2844 3798 2871 3816
rect 3096 3708 3123 3726
rect 3879 3843 3897 3870
rect 6093 3870 6120 3888
rect 6201 3870 6219 3888
rect 6093 3447 6111 3492
rect 1755 -1926 1773 -1899
rect 1728 -2133 1773 -2106
rect 3096 2646 3114 2682
rect 3051 2628 3069 2646
rect 3123 2529 3141 2547
rect 4491 3033 4518 3060
rect 3861 2997 3879 3024
rect 6183 3033 6201 3087
rect 3798 1701 3825 1728
rect 3096 1350 3114 1395
rect 2277 1017 2304 1035
rect 2241 936 2286 954
rect 3249 1008 3267 1044
rect 3096 324 3114 342
rect 2124 0 2160 18
rect 3888 324 3915 351
rect 3096 -621 3123 -603
rect 2079 -954 2097 -936
rect 1872 -3330 1890 -3285
rect 2196 -891 2214 -864
rect 2160 -2133 2178 -2106
rect 3879 -486 3897 -459
rect 6093 -459 6120 -441
rect 6201 -459 6219 -441
rect 6093 -882 6111 -837
rect 3096 -1683 3114 -1647
rect 3051 -1701 3069 -1683
rect 2799 -1764 2817 -1728
rect 3096 -1800 3114 -1764
rect 4491 -1296 4518 -1269
rect 3861 -1332 3879 -1305
rect 6183 -1296 6201 -1242
rect 3798 -2628 3825 -2601
rect 3096 -2979 3114 -2934
rect 2853 -4428 2871 -4401
rect 2196 -4761 2259 -4743
rect 2079 -5715 2097 -5697
rect 2853 -5373 2871 -5346
rect 2844 -7641 2871 -7623
<< metal2 >>
rect 1755 4743 2844 4761
rect 1755 18 1773 4743
rect 2196 63 2214 4572
rect 3096 4509 3114 4653
rect 3636 4653 3888 4680
rect 3636 4509 3654 4653
rect 3096 4491 3654 4509
rect 3771 3843 3879 3870
rect 2367 3798 2844 3816
rect 3105 3573 3123 3708
rect 3771 3573 3789 3843
rect 3105 3555 3789 3573
rect 6093 3492 6111 3870
rect 6183 3087 6201 3888
rect 3762 2997 3861 3024
rect 3051 2547 3069 2628
rect 3096 2547 3114 2646
rect 3762 2547 3780 2997
rect 3042 2511 3078 2547
rect 3096 2529 3123 2547
rect 3141 2529 3780 2547
rect 3051 2412 3069 2511
rect 4473 2412 4491 3060
rect 3051 2394 4491 2412
rect 3708 1701 3798 1728
rect 3096 1251 3114 1350
rect 3708 1251 3726 1701
rect 3096 1233 3726 1251
rect 3141 1035 3159 1233
rect 2304 1017 3159 1035
rect 3249 954 3267 1008
rect 2286 936 3267 954
rect 3096 180 3114 324
rect 3636 324 3888 351
rect 3636 180 3654 324
rect 3096 162 3654 180
rect 3096 63 3114 162
rect 2196 45 3114 63
rect 1755 0 2124 18
rect 1755 -1899 1773 0
rect 2196 -864 2214 45
rect 3771 -486 3879 -459
rect 3105 -756 3123 -621
rect 3771 -756 3789 -486
rect 3105 -774 3789 -756
rect 3105 -936 3123 -774
rect 6093 -837 6111 -459
rect 2097 -954 3123 -936
rect 6183 -1242 6201 -441
rect 3762 -1332 3861 -1305
rect 2799 -2106 2817 -1764
rect 3051 -1782 3069 -1701
rect 3096 -1764 3114 -1683
rect 3042 -1818 3078 -1782
rect 3762 -1782 3780 -1332
rect 3114 -1800 3780 -1782
rect 3051 -1917 3069 -1818
rect 4473 -1917 4491 -1269
rect 3051 -1935 4491 -1917
rect 1773 -2133 2160 -2106
rect 2178 -2133 2817 -2106
rect 3708 -2628 3798 -2601
rect 3096 -3078 3114 -2979
rect 3708 -3078 3726 -2628
rect 3096 -3096 3726 -3078
rect 3708 -3321 3726 -3096
rect 1890 -3330 3726 -3321
rect 1872 -3339 3726 -3330
rect 1872 -7623 1890 -3339
rect 2853 -4743 2871 -4428
rect 2259 -4761 2871 -4743
rect 2853 -5697 2871 -5373
rect 2097 -5715 2871 -5697
rect 1872 -7641 2844 -7623
<< m123contact >>
rect 3663 4968 3681 4995
rect 2403 4302 2421 4347
rect 2574 4329 2610 4347
rect 5157 4248 5175 4293
rect 3654 4023 3681 4050
rect 3627 3006 3654 3033
rect 4635 3033 4662 3060
rect 4896 3033 4923 3060
rect 2223 2340 2250 2358
rect 2313 2268 2331 2295
rect 2556 2277 2610 2295
rect 4338 1737 4365 1764
rect 4482 1737 4509 1764
rect 4608 1737 4635 1764
rect 4743 1737 4770 1764
rect 3051 1332 3069 1359
rect 3249 1053 3267 1071
rect 2223 1017 2250 1035
rect 3663 639 3681 666
rect 5157 -81 5175 -36
rect 3654 -306 3681 -279
rect 3627 -1323 3654 -1296
rect 4635 -1296 4662 -1269
rect 4896 -1296 4923 -1269
rect 1602 -2133 1620 -2106
rect 4338 -2592 4365 -2565
rect 4482 -2592 4509 -2565
rect 4608 -2592 4635 -2565
rect 4743 -2592 4770 -2565
rect 3051 -2997 3069 -2970
rect 1755 -4806 1773 -4788
rect 1809 -5751 1827 -5733
rect 3258 -4806 3276 -4788
rect 3258 -5751 3276 -5733
rect 1665 -7983 1683 -7938
<< metal3 >>
rect 2511 5310 3780 5328
rect 1602 2340 2223 2358
rect 1602 -2106 1620 2340
rect 1665 1017 2223 1035
rect 1665 -3258 1683 1017
rect 2313 -2052 2331 2268
rect 2403 -891 2421 4302
rect 2511 990 2529 5310
rect 3663 4950 3681 4968
rect 3762 4950 3780 5310
rect 3663 4932 3780 4950
rect 2610 4329 3456 4347
rect 3438 4266 3456 4329
rect 3663 4311 3681 4932
rect 3663 4293 5175 4311
rect 3438 4248 3771 4266
rect 3663 3996 3681 4023
rect 3753 3996 3771 4248
rect 3663 3978 3771 3996
rect 3663 3510 3681 3978
rect 3663 3492 4617 3510
rect 4599 3060 4617 3492
rect 4923 3339 4941 4293
rect 4851 3321 4941 3339
rect 4851 3060 4869 3321
rect 4599 3033 4635 3060
rect 4851 3033 4896 3060
rect 3654 3006 3690 3033
rect 3672 2295 3690 3006
rect 2610 2277 3690 2295
rect 3672 2079 3690 2277
rect 4599 2079 4617 3033
rect 3672 2061 4302 2079
rect 4284 1764 4302 2061
rect 4428 2061 4617 2079
rect 4428 1764 4446 2061
rect 4851 2034 4869 3033
rect 4581 2016 4869 2034
rect 4581 1764 4599 2016
rect 4284 1737 4338 1764
rect 4428 1737 4482 1764
rect 4581 1737 4608 1764
rect 4698 1737 4743 1764
rect 3051 1071 3069 1332
rect 4698 1071 4716 1737
rect 3051 1053 3249 1071
rect 3267 1053 4716 1071
rect 2511 972 3681 990
rect 3663 666 3681 972
rect 3663 -18 3681 639
rect 3663 -36 5175 -18
rect 3663 -819 3681 -306
rect 3663 -837 4617 -819
rect 3663 -891 3681 -837
rect 2403 -909 3681 -891
rect 4599 -1269 4617 -837
rect 4923 -990 4941 -36
rect 4851 -1008 4941 -990
rect 4851 -1269 4869 -1008
rect 4599 -1296 4635 -1269
rect 4851 -1296 4896 -1269
rect 3654 -1323 3690 -1296
rect 3672 -2052 3690 -1323
rect 2313 -2070 3690 -2052
rect 3672 -2250 3690 -2070
rect 4599 -2250 4617 -1296
rect 3672 -2268 4302 -2250
rect 4284 -2565 4302 -2268
rect 4428 -2268 4617 -2250
rect 4428 -2565 4446 -2268
rect 4851 -2295 4869 -1296
rect 4581 -2313 4869 -2295
rect 4581 -2565 4599 -2313
rect 4284 -2592 4338 -2565
rect 4428 -2592 4482 -2565
rect 4581 -2592 4608 -2565
rect 4698 -2592 4743 -2565
rect 3051 -3258 3069 -2997
rect 4698 -3258 4716 -2592
rect 1665 -3276 1755 -3258
rect 1773 -3276 4716 -3258
rect 1665 -7938 1683 -3276
rect 1773 -4806 3258 -4788
rect 1827 -5751 3258 -5733
<< labels >>
rlabel metal1 3168 1152 3168 1152 1 gnd
rlabel metal1 3447 1872 3447 1872 1 vdd
rlabel metal1 3645 1728 3645 1728 1 x0
rlabel m123contact 3636 3024 3636 3024 1 x1
rlabel metal1 3645 4041 3645 4041 1 x2
rlabel metal1 3636 4986 3636 4986 1 x3
rlabel polysilicon 3060 4761 3060 4761 1 a3
rlabel polysilicon 3060 4617 3060 4617 1 b3
rlabel metal1 3987 4671 3987 4671 1 a3_not
rlabel metal1 4824 4716 4824 4716 1 AlessB_3
rlabel polysilicon 3060 3681 3060 3681 1 b2
rlabel polysilicon 3060 3816 3060 3816 1 a2
rlabel metal1 3969 3870 3969 3870 1 a2_not
rlabel metal1 5580 3906 5580 3906 1 AlessB_2
rlabel metal1 6390 3852 6390 3852 7 AlessB
rlabel polysilicon 3060 2808 3060 2808 1 a1
rlabel polysilicon 3024 2628 3024 2628 1 b1
rlabel metal1 3951 3024 3951 3024 1 a1_not
rlabel metal1 5238 3078 5238 3078 1 AlessB_1
rlabel polysilicon 3051 1512 3051 1512 1 a0
rlabel polysilicon 3024 1332 3024 1332 1 b0
rlabel metal1 3906 1728 3906 1728 1 a0_not
rlabel metal1 5094 1782 5094 1782 1 AlessB_0
rlabel metal1 3987 351 3987 351 1 b3_not
rlabel metal1 3969 -459 3969 -459 1 b2_not
rlabel metal1 3951 -1305 3951 -1305 1 b1_not
rlabel metal1 3906 -2610 3906 -2610 1 b0_not
rlabel metal1 5085 -2538 5085 -2538 1 AmoreB_0
rlabel metal1 5256 -1251 5256 -1251 1 AmoreB_1
rlabel metal1 5589 -423 5589 -423 1 AmoreB_2
rlabel metal1 4833 378 4833 378 1 AmoreB_3
rlabel metal1 6399 -477 6399 -477 7 AmoreB
rlabel metal1 4770 -1287 4770 -1287 1 temp_more
rlabel metal1 4770 3042 4770 3042 1 temp_less
rlabel polycontact 5742 -5202 5742 -5202 1 k
rlabel polysilicon 5409 -5238 5409 -5238 1 temp
rlabel polysilicon 6381 -5220 6381 -5220 1 D2
rlabel metal1 6732 -5148 6732 -5148 1 AequalsB
rlabel m123contact 3669 -295 3669 -295 1 ab2xn
rlabel m123contact 3638 -1311 3644 -1308 1 ab1xn
rlabel m123contact 3672 652 3672 652 1 ab3xn
rlabel metal2 3854 -477 3854 -477 1 bh2
<< end >>
