magic
tech scmos
magscale 9 1
timestamp 1700484452
<< nwell >>
rect -92 15 -80 90
rect -53 85 -32 87
rect -53 83 -28 85
rect -53 82 -32 83
rect -52 70 -35 82
rect -52 69 -45 70
rect -43 69 -35 70
rect -92 -90 -80 -15
rect -53 -23 -32 -18
rect -52 -35 -35 -23
rect -52 -36 -45 -35
rect -43 -36 -35 -35
rect -92 -203 -80 -128
rect -53 -133 -32 -131
rect -30 -133 -28 -21
rect -53 -135 -28 -133
rect -53 -136 -32 -135
rect -52 -148 -35 -136
rect -52 -149 -45 -148
rect -43 -149 -35 -148
rect -92 -347 -80 -272
rect -53 -277 -32 -275
rect -30 -277 -28 -135
rect -53 -279 -28 -277
rect -53 -280 -32 -279
rect -52 -292 -35 -280
rect -52 -293 -45 -292
rect -43 -293 -35 -292
<< ntransistor >>
rect -117 81 -111 83
rect -117 62 -111 64
rect -45 60 -43 63
rect -117 40 -111 42
rect -117 22 -111 24
rect -117 -24 -111 -22
rect -117 -43 -111 -41
rect -45 -45 -43 -42
rect -117 -65 -111 -63
rect -117 -83 -111 -81
rect -117 -137 -111 -135
rect -117 -156 -111 -154
rect -45 -158 -43 -155
rect -117 -178 -111 -176
rect -117 -196 -111 -194
rect -117 -281 -111 -279
rect -117 -300 -111 -298
rect -45 -302 -43 -299
rect -117 -322 -111 -320
rect -117 -340 -111 -338
<< ptransistor >>
rect -89 81 -82 83
rect -45 71 -43 77
rect -89 62 -82 64
rect -89 40 -82 42
rect -89 22 -82 24
rect -89 -24 -82 -22
rect -45 -34 -43 -28
rect -89 -43 -82 -41
rect -89 -65 -82 -63
rect -89 -83 -82 -81
rect -89 -137 -82 -135
rect -45 -147 -43 -141
rect -89 -156 -82 -154
rect -89 -178 -82 -176
rect -89 -196 -82 -194
rect -89 -281 -82 -279
rect -45 -291 -43 -285
rect -89 -300 -82 -298
rect -89 -322 -82 -320
rect -89 -340 -82 -338
<< ndiffusion >>
rect -117 88 -111 89
rect -117 84 -116 88
rect -112 84 -111 88
rect -117 83 -111 84
rect -117 80 -111 81
rect -117 76 -116 80
rect -112 76 -111 80
rect -117 75 -111 76
rect -117 69 -111 70
rect -117 65 -116 69
rect -112 65 -111 69
rect -117 64 -111 65
rect -50 62 -45 63
rect -117 61 -111 62
rect -117 57 -116 61
rect -112 57 -111 61
rect -117 56 -111 57
rect -50 60 -49 62
rect -46 60 -45 62
rect -43 60 -41 63
rect -38 60 -37 63
rect -117 48 -111 49
rect -117 44 -116 48
rect -112 44 -111 48
rect -117 42 -111 44
rect -117 39 -111 40
rect -117 35 -116 39
rect -112 35 -111 39
rect -117 34 -111 35
rect -117 30 -111 31
rect -117 26 -116 30
rect -112 26 -111 30
rect -117 24 -111 26
rect -117 21 -111 22
rect -117 17 -116 21
rect -112 17 -111 21
rect -117 16 -111 17
rect -117 -17 -111 -16
rect -117 -21 -116 -17
rect -112 -21 -111 -17
rect -117 -22 -111 -21
rect -117 -25 -111 -24
rect -117 -29 -116 -25
rect -112 -29 -111 -25
rect -117 -30 -111 -29
rect -117 -36 -111 -35
rect -117 -40 -116 -36
rect -112 -40 -111 -36
rect -117 -41 -111 -40
rect -50 -43 -45 -42
rect -117 -44 -111 -43
rect -117 -48 -116 -44
rect -112 -48 -111 -44
rect -117 -49 -111 -48
rect -50 -45 -49 -43
rect -46 -45 -45 -43
rect -43 -45 -41 -42
rect -38 -45 -37 -42
rect -117 -57 -111 -56
rect -117 -61 -116 -57
rect -112 -61 -111 -57
rect -117 -63 -111 -61
rect -117 -66 -111 -65
rect -117 -70 -116 -66
rect -112 -70 -111 -66
rect -117 -71 -111 -70
rect -117 -75 -111 -74
rect -117 -79 -116 -75
rect -112 -79 -111 -75
rect -117 -81 -111 -79
rect -117 -84 -111 -83
rect -117 -88 -116 -84
rect -112 -88 -111 -84
rect -117 -89 -111 -88
rect -117 -130 -111 -129
rect -117 -134 -116 -130
rect -112 -134 -111 -130
rect -117 -135 -111 -134
rect -117 -138 -111 -137
rect -117 -142 -116 -138
rect -112 -142 -111 -138
rect -117 -143 -111 -142
rect -117 -149 -111 -148
rect -117 -153 -116 -149
rect -112 -153 -111 -149
rect -117 -154 -111 -153
rect -50 -156 -45 -155
rect -117 -157 -111 -156
rect -117 -161 -116 -157
rect -112 -161 -111 -157
rect -117 -162 -111 -161
rect -50 -158 -49 -156
rect -46 -158 -45 -156
rect -43 -158 -41 -155
rect -38 -158 -37 -155
rect -117 -170 -111 -169
rect -117 -174 -116 -170
rect -112 -174 -111 -170
rect -117 -176 -111 -174
rect -117 -179 -111 -178
rect -117 -183 -116 -179
rect -112 -183 -111 -179
rect -117 -184 -111 -183
rect -117 -188 -111 -187
rect -117 -192 -116 -188
rect -112 -192 -111 -188
rect -117 -194 -111 -192
rect -117 -197 -111 -196
rect -117 -201 -116 -197
rect -112 -201 -111 -197
rect -117 -202 -111 -201
rect -117 -274 -111 -273
rect -117 -278 -116 -274
rect -112 -278 -111 -274
rect -117 -279 -111 -278
rect -117 -282 -111 -281
rect -117 -286 -116 -282
rect -112 -286 -111 -282
rect -117 -287 -111 -286
rect -117 -293 -111 -292
rect -117 -297 -116 -293
rect -112 -297 -111 -293
rect -117 -298 -111 -297
rect -50 -300 -45 -299
rect -117 -301 -111 -300
rect -117 -305 -116 -301
rect -112 -305 -111 -301
rect -117 -306 -111 -305
rect -50 -302 -49 -300
rect -46 -302 -45 -300
rect -43 -302 -41 -299
rect -38 -302 -37 -299
rect -117 -314 -111 -313
rect -117 -318 -116 -314
rect -112 -318 -111 -314
rect -117 -320 -111 -318
rect -117 -323 -111 -322
rect -117 -327 -116 -323
rect -112 -327 -111 -323
rect -117 -328 -111 -327
rect -117 -332 -111 -331
rect -117 -336 -116 -332
rect -112 -336 -111 -332
rect -117 -338 -111 -336
rect -117 -341 -111 -340
rect -117 -345 -116 -341
rect -112 -345 -111 -341
rect -117 -346 -111 -345
<< pdiffusion >>
rect -89 88 -82 89
rect -89 84 -88 88
rect -84 84 -82 88
rect -89 83 -82 84
rect -89 80 -82 81
rect -89 76 -88 80
rect -84 76 -82 80
rect -89 75 -82 76
rect -89 69 -82 70
rect -89 65 -88 69
rect -84 65 -82 69
rect -89 64 -82 65
rect -50 74 -49 77
rect -46 74 -45 77
rect -50 71 -45 74
rect -43 76 -37 77
rect -43 73 -41 76
rect -38 73 -37 76
rect -43 71 -37 73
rect -89 61 -82 62
rect -89 57 -88 61
rect -84 57 -82 61
rect -89 56 -82 57
rect -89 48 -82 49
rect -89 44 -88 48
rect -84 44 -82 48
rect -89 42 -82 44
rect -89 39 -82 40
rect -89 35 -88 39
rect -84 35 -82 39
rect -89 34 -82 35
rect -89 30 -82 31
rect -89 26 -88 30
rect -84 26 -82 30
rect -89 24 -82 26
rect -89 21 -82 22
rect -89 17 -88 21
rect -84 17 -82 21
rect -89 16 -82 17
rect -89 -17 -82 -16
rect -89 -21 -88 -17
rect -84 -21 -82 -17
rect -89 -22 -82 -21
rect -89 -25 -82 -24
rect -89 -29 -88 -25
rect -84 -29 -82 -25
rect -89 -30 -82 -29
rect -89 -36 -82 -35
rect -89 -40 -88 -36
rect -84 -40 -82 -36
rect -89 -41 -82 -40
rect -50 -31 -49 -28
rect -46 -31 -45 -28
rect -50 -34 -45 -31
rect -43 -29 -37 -28
rect -43 -32 -41 -29
rect -38 -32 -37 -29
rect -43 -34 -37 -32
rect -89 -44 -82 -43
rect -89 -48 -88 -44
rect -84 -48 -82 -44
rect -89 -49 -82 -48
rect -89 -57 -82 -56
rect -89 -61 -88 -57
rect -84 -61 -82 -57
rect -89 -63 -82 -61
rect -89 -66 -82 -65
rect -89 -70 -88 -66
rect -84 -70 -82 -66
rect -89 -71 -82 -70
rect -89 -75 -82 -74
rect -89 -79 -88 -75
rect -84 -79 -82 -75
rect -89 -81 -82 -79
rect -89 -84 -82 -83
rect -89 -88 -88 -84
rect -84 -88 -82 -84
rect -89 -89 -82 -88
rect -89 -130 -82 -129
rect -89 -134 -88 -130
rect -84 -134 -82 -130
rect -89 -135 -82 -134
rect -89 -138 -82 -137
rect -89 -142 -88 -138
rect -84 -142 -82 -138
rect -89 -143 -82 -142
rect -89 -149 -82 -148
rect -89 -153 -88 -149
rect -84 -153 -82 -149
rect -89 -154 -82 -153
rect -50 -144 -49 -141
rect -46 -144 -45 -141
rect -50 -147 -45 -144
rect -43 -142 -37 -141
rect -43 -145 -41 -142
rect -38 -145 -37 -142
rect -43 -147 -37 -145
rect -89 -157 -82 -156
rect -89 -161 -88 -157
rect -84 -161 -82 -157
rect -89 -162 -82 -161
rect -89 -170 -82 -169
rect -89 -174 -88 -170
rect -84 -174 -82 -170
rect -89 -176 -82 -174
rect -89 -179 -82 -178
rect -89 -183 -88 -179
rect -84 -183 -82 -179
rect -89 -184 -82 -183
rect -89 -188 -82 -187
rect -89 -192 -88 -188
rect -84 -192 -82 -188
rect -89 -194 -82 -192
rect -89 -197 -82 -196
rect -89 -201 -88 -197
rect -84 -201 -82 -197
rect -89 -202 -82 -201
rect -89 -274 -82 -273
rect -89 -278 -88 -274
rect -84 -278 -82 -274
rect -89 -279 -82 -278
rect -89 -282 -82 -281
rect -89 -286 -88 -282
rect -84 -286 -82 -282
rect -89 -287 -82 -286
rect -89 -293 -82 -292
rect -89 -297 -88 -293
rect -84 -297 -82 -293
rect -89 -298 -82 -297
rect -50 -288 -49 -285
rect -46 -288 -45 -285
rect -50 -291 -45 -288
rect -43 -286 -37 -285
rect -43 -289 -41 -286
rect -38 -289 -37 -286
rect -43 -291 -37 -289
rect -89 -301 -82 -300
rect -89 -305 -88 -301
rect -84 -305 -82 -301
rect -89 -306 -82 -305
rect -89 -314 -82 -313
rect -89 -318 -88 -314
rect -84 -318 -82 -314
rect -89 -320 -82 -318
rect -89 -323 -82 -322
rect -89 -327 -88 -323
rect -84 -327 -82 -323
rect -89 -328 -82 -327
rect -89 -332 -82 -331
rect -89 -336 -88 -332
rect -84 -336 -82 -332
rect -89 -338 -82 -336
rect -89 -341 -82 -340
rect -89 -345 -88 -341
rect -84 -345 -82 -341
rect -89 -346 -82 -345
<< ndcontact >>
rect -116 84 -112 88
rect -116 76 -112 80
rect -116 65 -112 69
rect -116 57 -112 61
rect -49 59 -46 62
rect -41 60 -38 63
rect -116 44 -112 48
rect -116 35 -112 39
rect -116 26 -112 30
rect -116 17 -112 21
rect -116 -21 -112 -17
rect -116 -29 -112 -25
rect -116 -40 -112 -36
rect -116 -48 -112 -44
rect -49 -46 -46 -43
rect -41 -45 -38 -42
rect -116 -61 -112 -57
rect -116 -70 -112 -66
rect -116 -79 -112 -75
rect -116 -88 -112 -84
rect -116 -134 -112 -130
rect -116 -142 -112 -138
rect -116 -153 -112 -149
rect -116 -161 -112 -157
rect -49 -159 -46 -156
rect -41 -158 -38 -155
rect -116 -174 -112 -170
rect -116 -183 -112 -179
rect -116 -192 -112 -188
rect -116 -201 -112 -197
rect -116 -278 -112 -274
rect -116 -286 -112 -282
rect -116 -297 -112 -293
rect -116 -305 -112 -301
rect -49 -303 -46 -300
rect -41 -302 -38 -299
rect -116 -318 -112 -314
rect -116 -327 -112 -323
rect -116 -336 -112 -332
rect -116 -345 -112 -341
<< pdcontact >>
rect -88 84 -84 88
rect -88 76 -84 80
rect -88 65 -84 69
rect -49 74 -46 77
rect -41 73 -38 76
rect -88 57 -84 61
rect -88 44 -84 48
rect -88 35 -84 39
rect -88 26 -84 30
rect -88 17 -84 21
rect -88 -21 -84 -17
rect -88 -29 -84 -25
rect -88 -40 -84 -36
rect -49 -31 -46 -28
rect -41 -32 -38 -29
rect -88 -48 -84 -44
rect -88 -61 -84 -57
rect -88 -70 -84 -66
rect -88 -79 -84 -75
rect -88 -88 -84 -84
rect -88 -134 -84 -130
rect -88 -142 -84 -138
rect -88 -153 -84 -149
rect -49 -144 -46 -141
rect -41 -145 -38 -142
rect -88 -161 -84 -157
rect -88 -174 -84 -170
rect -88 -183 -84 -179
rect -88 -192 -84 -188
rect -88 -201 -84 -197
rect -88 -278 -84 -274
rect -88 -286 -84 -282
rect -88 -297 -84 -293
rect -49 -288 -46 -285
rect -41 -289 -38 -286
rect -88 -305 -84 -301
rect -88 -318 -84 -314
rect -88 -327 -84 -323
rect -88 -336 -84 -332
rect -88 -345 -84 -341
<< psubstratepcontact >>
rect -130 40 -126 44
rect -130 30 -126 34
rect -130 -65 -126 -61
rect -130 -75 -126 -71
rect -130 -178 -126 -174
rect -130 -188 -126 -184
rect -130 -322 -126 -318
rect -130 -332 -126 -328
<< nsubstratencontact >>
rect -75 40 -71 44
rect -75 30 -71 34
rect -75 -65 -71 -61
rect -75 -75 -71 -71
rect -75 -178 -71 -174
rect -75 -188 -71 -184
rect -75 -322 -71 -318
rect -75 -332 -71 -328
<< polysilicon >>
rect -123 93 -74 95
rect -123 83 -121 93
rect -140 81 -117 83
rect -111 81 -110 83
rect -108 81 -89 83
rect -82 81 -79 83
rect -140 10 -138 81
rect -108 64 -106 81
rect -76 64 -74 93
rect -45 77 -43 79
rect -45 67 -43 71
rect -135 62 -117 64
rect -111 62 -106 64
rect -93 62 -89 64
rect -82 62 -74 64
rect -69 64 -49 67
rect -44 64 -43 67
rect -45 63 -43 64
rect -135 24 -133 62
rect -45 58 -43 60
rect -103 42 -99 45
rect -124 40 -117 42
rect -111 40 -89 42
rect -82 40 -77 42
rect -103 24 -99 29
rect -135 22 -117 24
rect -111 22 -89 24
rect -82 22 -77 24
rect -140 8 -99 10
rect -123 -12 -74 -10
rect -123 -22 -121 -12
rect -140 -24 -117 -22
rect -111 -24 -110 -22
rect -108 -24 -89 -22
rect -82 -24 -79 -22
rect -140 -95 -138 -24
rect -108 -41 -106 -24
rect -76 -41 -74 -12
rect -45 -28 -43 -26
rect -45 -38 -43 -34
rect -135 -43 -117 -41
rect -111 -43 -106 -41
rect -93 -43 -89 -41
rect -82 -43 -74 -41
rect -69 -41 -49 -38
rect -44 -41 -43 -38
rect -45 -42 -43 -41
rect -135 -81 -133 -43
rect -45 -47 -43 -45
rect -103 -63 -99 -60
rect -124 -65 -117 -63
rect -111 -65 -89 -63
rect -82 -65 -77 -63
rect -103 -81 -99 -76
rect -135 -83 -117 -81
rect -111 -83 -89 -81
rect -82 -83 -77 -81
rect -140 -97 -99 -95
rect -123 -125 -74 -123
rect -123 -135 -121 -125
rect -140 -137 -117 -135
rect -111 -137 -110 -135
rect -108 -137 -89 -135
rect -82 -137 -79 -135
rect -140 -208 -138 -137
rect -108 -154 -106 -137
rect -76 -154 -74 -125
rect -45 -141 -43 -139
rect -45 -151 -43 -147
rect -135 -156 -117 -154
rect -111 -156 -106 -154
rect -93 -156 -89 -154
rect -82 -156 -74 -154
rect -69 -154 -49 -151
rect -44 -154 -43 -151
rect -45 -155 -43 -154
rect -135 -194 -133 -156
rect -45 -160 -43 -158
rect -103 -176 -99 -173
rect -124 -178 -117 -176
rect -111 -178 -89 -176
rect -82 -178 -77 -176
rect -103 -194 -99 -189
rect -135 -196 -117 -194
rect -111 -196 -89 -194
rect -82 -196 -77 -194
rect -140 -210 -99 -208
rect -123 -269 -74 -267
rect -123 -279 -121 -269
rect -140 -281 -117 -279
rect -111 -281 -110 -279
rect -108 -281 -89 -279
rect -82 -281 -79 -279
rect -140 -352 -138 -281
rect -108 -298 -106 -281
rect -76 -298 -74 -269
rect -45 -285 -43 -283
rect -45 -295 -43 -291
rect -135 -300 -117 -298
rect -111 -300 -106 -298
rect -93 -300 -89 -298
rect -82 -300 -74 -298
rect -69 -298 -49 -295
rect -44 -298 -43 -295
rect -45 -299 -43 -298
rect -135 -338 -133 -300
rect -45 -304 -43 -302
rect -103 -320 -99 -317
rect -124 -322 -117 -320
rect -111 -322 -89 -320
rect -82 -322 -77 -320
rect -103 -338 -99 -333
rect -135 -340 -117 -338
rect -111 -340 -89 -338
rect -82 -340 -77 -338
rect -140 -354 -99 -352
<< polycontact >>
rect -72 63 -69 67
rect -49 64 -44 67
rect -103 45 -99 49
rect -103 10 -99 14
rect -72 -42 -69 -38
rect -49 -41 -44 -38
rect -103 -60 -99 -56
rect -103 -95 -99 -91
rect -72 -155 -69 -151
rect -49 -154 -44 -151
rect -103 -173 -99 -169
rect -103 -208 -99 -204
rect -72 -299 -69 -295
rect -49 -298 -44 -295
rect -103 -317 -99 -313
rect -103 -352 -99 -348
<< metal1 >>
rect -112 84 -88 88
rect -84 84 -64 88
rect -112 76 -88 80
rect -84 76 -69 80
rect -130 65 -116 69
rect -112 65 -88 69
rect -73 67 -69 76
rect -130 54 -126 65
rect -73 63 -72 67
rect -73 61 -69 63
rect -112 57 -88 61
rect -84 57 -69 61
rect -68 54 -64 84
rect -130 50 -105 54
rect -130 44 -116 48
rect -130 38 -126 40
rect -109 39 -105 50
rect -103 50 -64 54
rect -60 83 -28 85
rect -103 49 -99 50
rect -84 44 -71 48
rect -148 36 -126 38
rect -148 4 -146 36
rect -130 34 -126 36
rect -112 35 -88 39
rect -75 38 -71 40
rect -60 38 -57 83
rect -50 82 -46 83
rect -49 77 -46 82
rect -41 68 -38 73
rect -41 65 -35 68
rect -41 63 -38 65
rect -49 56 -46 59
rect -75 35 -57 38
rect -52 54 -39 56
rect -75 34 -71 35
rect -130 26 -116 30
rect -84 26 -71 30
rect -112 17 -88 21
rect -103 14 -99 17
rect -52 4 -50 54
rect -148 2 -50 4
rect -148 -67 -146 2
rect -112 -21 -88 -17
rect -84 -21 -64 -17
rect -30 -20 -28 83
rect -112 -29 -88 -25
rect -84 -29 -69 -25
rect -130 -40 -116 -36
rect -112 -40 -88 -36
rect -73 -38 -69 -29
rect -130 -51 -126 -40
rect -73 -42 -72 -38
rect -73 -44 -69 -42
rect -112 -48 -88 -44
rect -84 -48 -69 -44
rect -68 -51 -64 -21
rect -130 -55 -105 -51
rect -130 -61 -116 -57
rect -130 -67 -126 -65
rect -109 -66 -105 -55
rect -103 -55 -64 -51
rect -60 -22 -28 -20
rect -103 -56 -99 -55
rect -84 -61 -71 -57
rect -148 -69 -126 -67
rect -148 -101 -146 -69
rect -130 -71 -126 -69
rect -112 -70 -88 -66
rect -75 -67 -71 -65
rect -60 -67 -57 -22
rect -50 -23 -46 -22
rect -49 -28 -46 -23
rect -41 -37 -38 -32
rect -41 -40 -35 -37
rect -41 -42 -38 -40
rect -49 -49 -46 -46
rect -75 -70 -57 -67
rect -52 -51 -39 -49
rect -75 -71 -71 -70
rect -130 -79 -116 -75
rect -84 -79 -71 -75
rect -112 -88 -88 -84
rect -103 -91 -99 -88
rect -52 -101 -50 -51
rect -148 -103 -50 -101
rect -148 -180 -146 -103
rect -112 -134 -88 -130
rect -84 -134 -64 -130
rect -30 -133 -28 -22
rect -112 -142 -88 -138
rect -84 -142 -69 -138
rect -130 -153 -116 -149
rect -112 -153 -88 -149
rect -73 -151 -69 -142
rect -130 -164 -126 -153
rect -73 -155 -72 -151
rect -73 -157 -69 -155
rect -112 -161 -88 -157
rect -84 -161 -69 -157
rect -68 -164 -64 -134
rect -130 -168 -105 -164
rect -130 -174 -116 -170
rect -130 -180 -126 -178
rect -109 -179 -105 -168
rect -103 -168 -64 -164
rect -60 -135 -28 -133
rect -103 -169 -99 -168
rect -84 -174 -71 -170
rect -148 -182 -126 -180
rect -148 -214 -146 -182
rect -130 -184 -126 -182
rect -112 -183 -88 -179
rect -75 -180 -71 -178
rect -60 -180 -57 -135
rect -50 -136 -46 -135
rect -49 -141 -46 -136
rect -41 -150 -38 -145
rect -41 -153 -35 -150
rect -41 -155 -38 -153
rect -49 -162 -46 -159
rect -75 -183 -57 -180
rect -52 -164 -39 -162
rect -75 -184 -71 -183
rect -130 -192 -116 -188
rect -84 -192 -71 -188
rect -112 -201 -88 -197
rect -103 -204 -99 -201
rect -52 -214 -50 -164
rect -148 -216 -50 -214
rect -148 -324 -146 -216
rect -112 -278 -88 -274
rect -84 -278 -64 -274
rect -30 -277 -28 -135
rect -112 -286 -88 -282
rect -84 -286 -69 -282
rect -130 -297 -116 -293
rect -112 -297 -88 -293
rect -73 -295 -69 -286
rect -130 -308 -126 -297
rect -73 -299 -72 -295
rect -73 -301 -69 -299
rect -112 -305 -88 -301
rect -84 -305 -69 -301
rect -68 -308 -64 -278
rect -130 -312 -105 -308
rect -130 -318 -116 -314
rect -130 -324 -126 -322
rect -109 -323 -105 -312
rect -103 -312 -64 -308
rect -60 -279 -28 -277
rect -103 -313 -99 -312
rect -84 -318 -71 -314
rect -148 -326 -126 -324
rect -148 -358 -146 -326
rect -130 -328 -126 -326
rect -112 -327 -88 -323
rect -75 -324 -71 -322
rect -60 -324 -57 -279
rect -50 -280 -46 -279
rect -49 -285 -46 -280
rect -41 -294 -38 -289
rect -41 -297 -35 -294
rect -41 -299 -38 -297
rect -49 -306 -46 -303
rect -75 -327 -57 -324
rect -52 -308 -39 -306
rect -75 -328 -71 -327
rect -130 -336 -116 -332
rect -84 -336 -71 -332
rect -112 -345 -88 -341
rect -103 -348 -99 -345
rect -52 -358 -50 -308
rect -148 -360 -50 -358
<< labels >>
rlabel metal1 -89 -359 -89 -359 1 gnd
rlabel metal1 -58 -279 -58 -279 1 vdd
rlabel metal1 -36 -295 -36 -295 1 x0
rlabel polysilicon -101 -320 -101 -320 1 b0
rlabel polysilicon -101 -338 -101 -338 1 a0
rlabel polysilicon -101 -193 -101 -193 1 a1
rlabel polysilicon -102 -176 -102 -176 1 b1
rlabel metal1 -37 -151 -37 -151 1 x1
rlabel polysilicon -101 -79 -101 -79 1 a2
rlabel polysilicon -101 -62 -101 -62 1 b2
rlabel metal1 -36 -38 -36 -38 1 x2
rlabel polysilicon -101 25 -101 25 1 a3
rlabel polysilicon -101 44 -101 44 1 b3
rlabel metal1 -37 67 -37 67 1 x3
<< end >>
