magic
tech scmos
magscale 9 1
timestamp 1700922445
<< nwell >>
rect -523 300 -511 375
rect -484 367 -463 372
rect -483 355 -466 367
rect -483 354 -476 355
rect -474 354 -466 355
rect -443 333 -422 338
rect -349 337 -328 343
rect -442 321 -425 333
rect -442 320 -435 321
rect -433 320 -425 321
rect -401 320 -365 330
rect -349 325 -332 337
rect -349 324 -342 325
rect -340 324 -332 325
rect -523 195 -511 270
rect -484 262 -463 267
rect -483 250 -466 262
rect -483 249 -476 250
rect -474 249 -466 250
rect -445 245 -424 248
rect -446 243 -424 245
rect -357 247 -336 253
rect -265 250 -244 253
rect -265 248 -213 250
rect -265 247 -244 248
rect -444 231 -427 243
rect -444 230 -437 231
rect -435 230 -427 231
rect -409 230 -373 240
rect -357 235 -340 247
rect -357 234 -350 235
rect -348 234 -340 235
rect -317 230 -281 240
rect -265 235 -248 247
rect -215 243 -213 248
rect -265 234 -258 235
rect -256 234 -248 235
rect -217 230 -159 243
rect -183 228 -179 230
rect -393 159 -283 162
rect -523 82 -511 157
rect -394 156 -283 159
rect -484 149 -464 154
rect -447 149 -426 154
rect -483 137 -466 149
rect -483 136 -476 137
rect -474 136 -466 137
rect -446 137 -429 149
rect -393 144 -283 156
rect -446 136 -439 137
rect -437 136 -429 137
rect -410 15 -300 18
rect -523 -62 -511 13
rect -411 12 -300 15
rect -484 5 -464 10
rect -453 5 -432 10
rect -483 -7 -466 5
rect -483 -8 -476 -7
rect -474 -8 -466 -7
rect -452 -7 -435 5
rect -410 0 -300 12
rect -452 -8 -445 -7
rect -443 -8 -435 -7
<< ntransistor >>
rect -548 366 -542 368
rect -548 347 -542 349
rect -476 345 -474 348
rect -548 325 -542 327
rect -548 307 -542 309
rect -435 311 -433 314
rect -342 315 -340 318
rect -393 309 -391 312
rect -381 309 -380 312
rect -375 309 -373 312
rect -548 261 -542 263
rect -548 242 -542 244
rect -476 240 -474 243
rect -548 220 -542 222
rect -437 221 -435 224
rect -350 225 -348 228
rect -258 225 -256 228
rect -401 219 -399 222
rect -389 219 -388 222
rect -383 219 -381 222
rect -309 219 -307 222
rect -291 219 -289 222
rect -211 219 -209 222
rect -201 219 -199 222
rect -191 219 -189 222
rect -181 219 -179 222
rect -167 219 -165 222
rect -548 202 -542 204
rect -548 148 -542 150
rect -548 129 -542 131
rect -476 127 -474 130
rect -439 127 -437 130
rect -383 129 -381 132
rect -369 129 -367 132
rect -353 129 -351 132
rect -339 129 -337 132
rect -324 129 -322 132
rect -295 129 -293 132
rect -548 107 -542 109
rect -548 89 -542 91
rect -548 4 -542 6
rect -548 -15 -542 -13
rect -476 -17 -474 -14
rect -445 -17 -443 -14
rect -400 -15 -398 -12
rect -386 -15 -384 -12
rect -370 -15 -368 -12
rect -356 -15 -354 -12
rect -341 -15 -339 -12
rect -312 -15 -310 -12
rect -548 -37 -542 -35
rect -548 -55 -542 -53
<< ptransistor >>
rect -520 366 -513 368
rect -476 356 -474 362
rect -520 347 -513 349
rect -520 325 -513 327
rect -520 307 -513 309
rect -435 322 -433 328
rect -393 323 -391 328
rect -375 323 -373 328
rect -342 326 -340 332
rect -520 261 -513 263
rect -476 251 -474 257
rect -520 242 -513 244
rect -520 220 -513 222
rect -437 232 -435 238
rect -401 233 -399 238
rect -383 233 -381 238
rect -350 236 -348 242
rect -309 233 -307 238
rect -291 233 -289 238
rect -258 236 -256 242
rect -211 232 -209 237
rect -205 232 -203 237
rect -201 232 -199 237
rect -191 232 -189 237
rect -181 232 -179 237
rect -167 232 -165 237
rect -520 202 -513 204
rect -520 148 -513 150
rect -383 146 -381 152
rect -369 146 -367 152
rect -353 146 -351 152
rect -339 146 -337 152
rect -324 146 -322 152
rect -295 146 -293 152
rect -476 138 -474 144
rect -439 138 -437 144
rect -520 129 -513 131
rect -520 107 -513 109
rect -520 89 -513 91
rect -520 4 -513 6
rect -400 2 -398 8
rect -386 2 -384 8
rect -370 2 -368 8
rect -356 2 -354 8
rect -341 2 -339 8
rect -312 2 -310 8
rect -476 -6 -474 0
rect -445 -6 -443 0
rect -520 -15 -513 -13
rect -520 -37 -513 -35
rect -520 -55 -513 -53
<< ndiffusion >>
rect -548 373 -542 374
rect -548 369 -547 373
rect -543 369 -542 373
rect -548 368 -542 369
rect -548 365 -542 366
rect -548 361 -547 365
rect -543 361 -542 365
rect -548 360 -542 361
rect -548 354 -542 355
rect -548 350 -547 354
rect -543 350 -542 354
rect -548 349 -542 350
rect -481 347 -476 348
rect -548 346 -542 347
rect -548 342 -547 346
rect -543 342 -542 346
rect -548 341 -542 342
rect -481 345 -480 347
rect -477 345 -476 347
rect -474 345 -472 348
rect -469 345 -468 348
rect -548 333 -542 334
rect -548 329 -547 333
rect -543 329 -542 333
rect -548 327 -542 329
rect -548 324 -542 325
rect -548 320 -547 324
rect -543 320 -542 324
rect -548 319 -542 320
rect -548 315 -542 316
rect -548 311 -547 315
rect -543 311 -542 315
rect -548 309 -542 311
rect -548 306 -542 307
rect -548 302 -547 306
rect -543 302 -542 306
rect -548 301 -542 302
rect -440 313 -435 314
rect -440 311 -439 313
rect -436 311 -435 313
rect -433 311 -431 314
rect -428 311 -427 314
rect -347 317 -342 318
rect -347 315 -346 317
rect -343 315 -342 317
rect -340 315 -338 318
rect -335 315 -334 318
rect -397 311 -393 312
rect -397 309 -396 311
rect -394 309 -393 311
rect -391 309 -381 312
rect -380 309 -375 312
rect -373 310 -372 312
rect -370 310 -369 312
rect -373 309 -369 310
rect -548 268 -542 269
rect -548 264 -547 268
rect -543 264 -542 268
rect -548 263 -542 264
rect -548 260 -542 261
rect -548 256 -547 260
rect -543 256 -542 260
rect -548 255 -542 256
rect -548 249 -542 250
rect -548 245 -547 249
rect -543 245 -542 249
rect -548 244 -542 245
rect -481 242 -476 243
rect -548 241 -542 242
rect -548 237 -547 241
rect -543 237 -542 241
rect -548 236 -542 237
rect -481 240 -480 242
rect -477 240 -476 242
rect -474 240 -472 243
rect -469 240 -468 243
rect -548 228 -542 229
rect -548 224 -547 228
rect -543 224 -542 228
rect -548 222 -542 224
rect -548 219 -542 220
rect -548 215 -547 219
rect -543 215 -542 219
rect -548 214 -542 215
rect -442 223 -437 224
rect -442 221 -441 223
rect -438 221 -437 223
rect -435 221 -433 224
rect -430 221 -429 224
rect -355 227 -350 228
rect -355 225 -354 227
rect -351 225 -350 227
rect -348 225 -346 228
rect -343 225 -342 228
rect -263 227 -258 228
rect -263 225 -262 227
rect -259 225 -258 227
rect -256 225 -254 228
rect -251 225 -250 228
rect -405 221 -401 222
rect -405 219 -404 221
rect -402 219 -401 221
rect -399 219 -389 222
rect -388 219 -383 222
rect -381 220 -380 222
rect -378 220 -377 222
rect -381 219 -377 220
rect -313 221 -309 222
rect -313 219 -312 221
rect -310 219 -309 221
rect -307 219 -291 222
rect -289 220 -288 222
rect -286 220 -285 222
rect -289 219 -285 220
rect -216 220 -215 222
rect -213 220 -211 222
rect -216 219 -211 220
rect -209 220 -208 222
rect -209 219 -206 220
rect -205 220 -204 222
rect -202 220 -201 222
rect -205 219 -201 220
rect -199 220 -198 222
rect -199 219 -196 220
rect -195 220 -194 222
rect -192 220 -191 222
rect -195 219 -191 220
rect -189 220 -188 222
rect -189 219 -186 220
rect -185 220 -184 222
rect -182 220 -181 222
rect -185 219 -181 220
rect -179 220 -178 222
rect -179 219 -176 220
rect -171 220 -170 222
rect -168 220 -167 222
rect -171 219 -167 220
rect -165 220 -164 222
rect -162 220 -161 222
rect -165 219 -161 220
rect -548 210 -542 211
rect -548 206 -547 210
rect -543 206 -542 210
rect -548 204 -542 206
rect -548 201 -542 202
rect -548 197 -547 201
rect -543 197 -542 201
rect -548 196 -542 197
rect -548 155 -542 156
rect -548 151 -547 155
rect -543 151 -542 155
rect -548 150 -542 151
rect -548 147 -542 148
rect -548 143 -547 147
rect -543 143 -542 147
rect -548 142 -542 143
rect -548 136 -542 137
rect -548 132 -547 136
rect -543 132 -542 136
rect -548 131 -542 132
rect -481 129 -476 130
rect -548 128 -542 129
rect -548 124 -547 128
rect -543 124 -542 128
rect -548 123 -542 124
rect -481 127 -480 129
rect -477 127 -476 129
rect -474 127 -472 130
rect -469 127 -468 130
rect -444 129 -439 130
rect -444 127 -443 129
rect -440 127 -439 129
rect -437 127 -435 130
rect -432 127 -431 130
rect -388 129 -387 132
rect -384 129 -383 132
rect -381 129 -369 132
rect -367 129 -353 132
rect -351 129 -339 132
rect -337 129 -324 132
rect -322 129 -318 132
rect -315 129 -307 132
rect -301 129 -299 132
rect -296 129 -295 132
rect -293 129 -292 132
rect -289 129 -288 132
rect -548 115 -542 116
rect -548 111 -547 115
rect -543 111 -542 115
rect -548 109 -542 111
rect -548 106 -542 107
rect -548 102 -547 106
rect -543 102 -542 106
rect -548 101 -542 102
rect -548 97 -542 98
rect -548 93 -547 97
rect -543 93 -542 97
rect -548 91 -542 93
rect -548 88 -542 89
rect -548 84 -547 88
rect -543 84 -542 88
rect -548 83 -542 84
rect -548 11 -542 12
rect -548 7 -547 11
rect -543 7 -542 11
rect -548 6 -542 7
rect -548 3 -542 4
rect -548 -1 -547 3
rect -543 -1 -542 3
rect -548 -2 -542 -1
rect -548 -8 -542 -7
rect -548 -12 -547 -8
rect -543 -12 -542 -8
rect -548 -13 -542 -12
rect -481 -15 -476 -14
rect -548 -16 -542 -15
rect -548 -20 -547 -16
rect -543 -20 -542 -16
rect -548 -21 -542 -20
rect -481 -17 -480 -15
rect -477 -17 -476 -15
rect -474 -17 -472 -14
rect -469 -17 -468 -14
rect -450 -15 -445 -14
rect -450 -17 -449 -15
rect -446 -17 -445 -15
rect -443 -17 -441 -14
rect -438 -17 -437 -14
rect -405 -15 -404 -12
rect -401 -15 -400 -12
rect -398 -15 -386 -12
rect -384 -15 -370 -12
rect -368 -15 -356 -12
rect -354 -15 -341 -12
rect -339 -15 -335 -12
rect -332 -15 -324 -12
rect -318 -15 -316 -12
rect -313 -15 -312 -12
rect -310 -15 -309 -12
rect -306 -15 -305 -12
rect -548 -29 -542 -28
rect -548 -33 -547 -29
rect -543 -33 -542 -29
rect -548 -35 -542 -33
rect -548 -38 -542 -37
rect -548 -42 -547 -38
rect -543 -42 -542 -38
rect -548 -43 -542 -42
rect -548 -47 -542 -46
rect -548 -51 -547 -47
rect -543 -51 -542 -47
rect -548 -53 -542 -51
rect -548 -56 -542 -55
rect -548 -60 -547 -56
rect -543 -60 -542 -56
rect -548 -61 -542 -60
<< pdiffusion >>
rect -520 373 -513 374
rect -520 369 -519 373
rect -515 369 -513 373
rect -520 368 -513 369
rect -520 365 -513 366
rect -520 361 -519 365
rect -515 361 -513 365
rect -520 360 -513 361
rect -520 354 -513 355
rect -520 350 -519 354
rect -515 350 -513 354
rect -520 349 -513 350
rect -481 359 -480 362
rect -477 359 -476 362
rect -481 356 -476 359
rect -474 361 -468 362
rect -474 358 -472 361
rect -469 358 -468 361
rect -474 356 -468 358
rect -520 346 -513 347
rect -520 342 -519 346
rect -515 342 -513 346
rect -520 341 -513 342
rect -520 333 -513 334
rect -520 329 -519 333
rect -515 329 -513 333
rect -520 327 -513 329
rect -520 324 -513 325
rect -520 320 -519 324
rect -515 320 -513 324
rect -520 319 -513 320
rect -520 315 -513 316
rect -520 311 -519 315
rect -515 311 -513 315
rect -520 309 -513 311
rect -520 306 -513 307
rect -520 302 -519 306
rect -515 302 -513 306
rect -520 301 -513 302
rect -347 329 -346 332
rect -343 329 -342 332
rect -440 325 -439 328
rect -436 325 -435 328
rect -440 322 -435 325
rect -433 327 -427 328
rect -433 324 -431 327
rect -428 324 -427 327
rect -433 322 -427 324
rect -397 327 -393 328
rect -397 325 -396 327
rect -394 325 -393 327
rect -397 323 -393 325
rect -391 326 -384 328
rect -391 324 -390 326
rect -388 324 -384 326
rect -391 323 -384 324
rect -380 327 -375 328
rect -380 325 -379 327
rect -377 325 -375 327
rect -380 323 -375 325
rect -373 327 -369 328
rect -373 325 -372 327
rect -370 325 -369 327
rect -347 326 -342 329
rect -340 331 -334 332
rect -340 328 -338 331
rect -335 328 -334 331
rect -340 326 -334 328
rect -373 323 -369 325
rect -520 268 -513 269
rect -520 264 -519 268
rect -515 264 -513 268
rect -520 263 -513 264
rect -520 260 -513 261
rect -520 256 -519 260
rect -515 256 -513 260
rect -520 255 -513 256
rect -520 249 -513 250
rect -520 245 -519 249
rect -515 245 -513 249
rect -520 244 -513 245
rect -481 254 -480 257
rect -477 254 -476 257
rect -481 251 -476 254
rect -474 256 -468 257
rect -474 253 -472 256
rect -469 253 -468 256
rect -474 251 -468 253
rect -520 241 -513 242
rect -520 237 -519 241
rect -515 237 -513 241
rect -355 239 -354 242
rect -351 239 -350 242
rect -520 236 -513 237
rect -520 228 -513 229
rect -520 224 -519 228
rect -515 224 -513 228
rect -520 222 -513 224
rect -520 219 -513 220
rect -520 215 -519 219
rect -515 215 -513 219
rect -442 235 -441 238
rect -438 235 -437 238
rect -442 232 -437 235
rect -435 237 -429 238
rect -435 234 -433 237
rect -430 234 -429 237
rect -435 232 -429 234
rect -405 237 -401 238
rect -405 235 -404 237
rect -402 235 -401 237
rect -405 233 -401 235
rect -399 236 -392 238
rect -399 234 -398 236
rect -396 234 -392 236
rect -399 233 -392 234
rect -388 237 -383 238
rect -388 235 -387 237
rect -385 235 -383 237
rect -388 233 -383 235
rect -381 237 -377 238
rect -381 235 -380 237
rect -378 235 -377 237
rect -355 236 -350 239
rect -348 241 -342 242
rect -348 238 -346 241
rect -343 238 -342 241
rect -348 236 -342 238
rect -313 237 -309 238
rect -381 233 -377 235
rect -313 235 -312 237
rect -310 235 -309 237
rect -313 233 -309 235
rect -307 236 -300 238
rect -307 234 -306 236
rect -304 234 -300 236
rect -307 233 -300 234
rect -263 239 -262 242
rect -259 239 -258 242
rect -296 237 -291 238
rect -296 235 -295 237
rect -293 235 -291 237
rect -296 233 -291 235
rect -289 237 -285 238
rect -289 235 -288 237
rect -286 235 -285 237
rect -263 236 -258 239
rect -256 241 -250 242
rect -256 238 -254 241
rect -251 238 -250 241
rect -256 236 -250 238
rect -216 236 -211 237
rect -289 233 -285 235
rect -216 234 -215 236
rect -213 234 -211 236
rect -216 232 -211 234
rect -209 232 -205 237
rect -203 232 -201 237
rect -199 232 -191 237
rect -189 232 -181 237
rect -179 235 -176 237
rect -179 233 -178 235
rect -179 232 -176 233
rect -171 236 -167 237
rect -171 234 -170 236
rect -168 234 -167 236
rect -171 232 -167 234
rect -165 235 -161 237
rect -165 233 -164 235
rect -162 233 -161 235
rect -165 232 -161 233
rect -520 214 -513 215
rect -520 210 -513 211
rect -520 206 -519 210
rect -515 206 -513 210
rect -520 204 -513 206
rect -520 201 -513 202
rect -520 197 -519 201
rect -515 197 -513 201
rect -520 196 -513 197
rect -520 155 -513 156
rect -520 151 -519 155
rect -515 151 -513 155
rect -520 150 -513 151
rect -520 147 -513 148
rect -520 143 -519 147
rect -515 143 -513 147
rect -520 142 -513 143
rect -520 136 -513 137
rect -520 132 -519 136
rect -515 132 -513 136
rect -520 131 -513 132
rect -388 151 -383 152
rect -388 148 -387 151
rect -384 148 -383 151
rect -388 146 -383 148
rect -381 150 -376 152
rect -381 147 -380 150
rect -377 147 -376 150
rect -381 146 -376 147
rect -374 151 -369 152
rect -374 148 -373 151
rect -370 148 -369 151
rect -374 146 -369 148
rect -367 150 -361 152
rect -367 147 -366 150
rect -363 147 -361 150
rect -367 146 -361 147
rect -359 151 -353 152
rect -359 148 -357 151
rect -354 148 -353 151
rect -359 146 -353 148
rect -351 150 -346 152
rect -351 147 -350 150
rect -347 147 -346 150
rect -351 146 -346 147
rect -344 151 -339 152
rect -344 148 -343 151
rect -340 148 -339 151
rect -344 146 -339 148
rect -337 150 -332 152
rect -337 147 -336 150
rect -333 147 -332 150
rect -337 146 -332 147
rect -330 151 -324 152
rect -330 148 -329 151
rect -326 148 -324 151
rect -330 146 -324 148
rect -322 150 -307 152
rect -322 147 -321 150
rect -318 147 -307 150
rect -322 146 -307 147
rect -301 149 -299 152
rect -296 149 -295 152
rect -301 146 -295 149
rect -293 150 -288 152
rect -293 147 -292 150
rect -289 147 -288 150
rect -293 146 -288 147
rect -481 141 -480 144
rect -477 141 -476 144
rect -481 138 -476 141
rect -474 143 -468 144
rect -474 140 -472 143
rect -469 140 -468 143
rect -474 138 -468 140
rect -444 141 -443 144
rect -440 141 -439 144
rect -444 138 -439 141
rect -437 143 -431 144
rect -437 140 -435 143
rect -432 140 -431 143
rect -437 138 -431 140
rect -520 128 -513 129
rect -520 124 -519 128
rect -515 124 -513 128
rect -520 123 -513 124
rect -520 115 -513 116
rect -520 111 -519 115
rect -515 111 -513 115
rect -520 109 -513 111
rect -520 106 -513 107
rect -520 102 -519 106
rect -515 102 -513 106
rect -520 101 -513 102
rect -520 97 -513 98
rect -520 93 -519 97
rect -515 93 -513 97
rect -520 91 -513 93
rect -520 88 -513 89
rect -520 84 -519 88
rect -515 84 -513 88
rect -520 83 -513 84
rect -520 11 -513 12
rect -520 7 -519 11
rect -515 7 -513 11
rect -520 6 -513 7
rect -520 3 -513 4
rect -520 -1 -519 3
rect -515 -1 -513 3
rect -520 -2 -513 -1
rect -520 -8 -513 -7
rect -520 -12 -519 -8
rect -515 -12 -513 -8
rect -520 -13 -513 -12
rect -405 7 -400 8
rect -405 4 -404 7
rect -401 4 -400 7
rect -405 2 -400 4
rect -398 6 -393 8
rect -398 3 -397 6
rect -394 3 -393 6
rect -398 2 -393 3
rect -391 7 -386 8
rect -391 4 -390 7
rect -387 4 -386 7
rect -391 2 -386 4
rect -384 6 -378 8
rect -384 3 -383 6
rect -380 3 -378 6
rect -384 2 -378 3
rect -376 7 -370 8
rect -376 4 -374 7
rect -371 4 -370 7
rect -376 2 -370 4
rect -368 6 -363 8
rect -368 3 -367 6
rect -364 3 -363 6
rect -368 2 -363 3
rect -361 7 -356 8
rect -361 4 -360 7
rect -357 4 -356 7
rect -361 2 -356 4
rect -354 6 -349 8
rect -354 3 -353 6
rect -350 3 -349 6
rect -354 2 -349 3
rect -347 7 -341 8
rect -347 4 -346 7
rect -343 4 -341 7
rect -347 2 -341 4
rect -339 6 -324 8
rect -339 3 -338 6
rect -335 3 -324 6
rect -339 2 -324 3
rect -318 5 -316 8
rect -313 5 -312 8
rect -318 2 -312 5
rect -310 6 -305 8
rect -310 3 -309 6
rect -306 3 -305 6
rect -310 2 -305 3
rect -481 -3 -480 0
rect -477 -3 -476 0
rect -481 -6 -476 -3
rect -474 -1 -468 0
rect -474 -4 -472 -1
rect -469 -4 -468 -1
rect -474 -6 -468 -4
rect -450 -3 -449 0
rect -446 -3 -445 0
rect -450 -6 -445 -3
rect -443 -1 -437 0
rect -443 -4 -441 -1
rect -438 -4 -437 -1
rect -443 -6 -437 -4
rect -520 -16 -513 -15
rect -520 -20 -519 -16
rect -515 -20 -513 -16
rect -520 -21 -513 -20
rect -520 -29 -513 -28
rect -520 -33 -519 -29
rect -515 -33 -513 -29
rect -520 -35 -513 -33
rect -520 -38 -513 -37
rect -520 -42 -519 -38
rect -515 -42 -513 -38
rect -520 -43 -513 -42
rect -520 -47 -513 -46
rect -520 -51 -519 -47
rect -515 -51 -513 -47
rect -520 -53 -513 -51
rect -520 -56 -513 -55
rect -520 -60 -519 -56
rect -515 -60 -513 -56
rect -520 -61 -513 -60
<< ndcontact >>
rect -547 369 -543 373
rect -547 361 -543 365
rect -547 350 -543 354
rect -547 342 -543 346
rect -480 344 -477 347
rect -472 345 -469 348
rect -547 329 -543 333
rect -547 320 -543 324
rect -547 311 -543 315
rect -547 302 -543 306
rect -439 310 -436 313
rect -431 311 -428 314
rect -346 314 -343 317
rect -338 315 -335 318
rect -396 309 -394 311
rect -372 310 -370 312
rect -547 264 -543 268
rect -547 256 -543 260
rect -547 245 -543 249
rect -547 237 -543 241
rect -480 239 -477 242
rect -472 240 -469 243
rect -547 224 -543 228
rect -547 215 -543 219
rect -441 220 -438 223
rect -433 221 -430 224
rect -354 224 -351 227
rect -346 225 -343 228
rect -262 224 -259 227
rect -254 225 -251 228
rect -404 219 -402 221
rect -380 220 -378 222
rect -312 219 -310 221
rect -288 220 -286 222
rect -215 220 -213 222
rect -208 220 -206 222
rect -204 220 -202 222
rect -198 220 -196 222
rect -194 220 -192 222
rect -188 220 -186 222
rect -184 220 -182 222
rect -178 220 -176 222
rect -170 220 -168 222
rect -164 220 -162 222
rect -547 206 -543 210
rect -547 197 -543 201
rect -547 151 -543 155
rect -547 143 -543 147
rect -547 132 -543 136
rect -547 124 -543 128
rect -480 126 -477 129
rect -472 127 -469 130
rect -443 126 -440 129
rect -435 127 -432 130
rect -387 129 -384 132
rect -318 129 -315 132
rect -299 129 -296 132
rect -292 129 -289 132
rect -547 111 -543 115
rect -547 102 -543 106
rect -547 93 -543 97
rect -547 84 -543 88
rect -547 7 -543 11
rect -547 -1 -543 3
rect -547 -12 -543 -8
rect -547 -20 -543 -16
rect -480 -18 -477 -15
rect -472 -17 -469 -14
rect -449 -18 -446 -15
rect -441 -17 -438 -14
rect -404 -15 -401 -12
rect -335 -15 -332 -12
rect -316 -15 -313 -12
rect -309 -15 -306 -12
rect -547 -33 -543 -29
rect -547 -42 -543 -38
rect -547 -51 -543 -47
rect -547 -60 -543 -56
<< pdcontact >>
rect -519 369 -515 373
rect -519 361 -515 365
rect -519 350 -515 354
rect -480 359 -477 362
rect -472 358 -469 361
rect -519 342 -515 346
rect -519 329 -515 333
rect -519 320 -515 324
rect -519 311 -515 315
rect -519 302 -515 306
rect -346 329 -343 332
rect -439 325 -436 328
rect -431 324 -428 327
rect -396 325 -394 327
rect -390 324 -388 326
rect -379 325 -377 327
rect -372 325 -370 327
rect -338 328 -335 331
rect -519 264 -515 268
rect -519 256 -515 260
rect -519 245 -515 249
rect -480 254 -477 257
rect -472 253 -469 256
rect -519 237 -515 241
rect -354 239 -351 242
rect -519 224 -515 228
rect -519 215 -515 219
rect -441 235 -438 238
rect -433 234 -430 237
rect -404 235 -402 237
rect -398 234 -396 236
rect -387 235 -385 237
rect -380 235 -378 237
rect -346 238 -343 241
rect -312 235 -310 237
rect -306 234 -304 236
rect -262 239 -259 242
rect -295 235 -293 237
rect -288 235 -286 237
rect -254 238 -251 241
rect -215 234 -213 236
rect -178 233 -176 235
rect -170 234 -168 236
rect -164 233 -162 235
rect -519 206 -515 210
rect -519 197 -515 201
rect -519 151 -515 155
rect -519 143 -515 147
rect -519 132 -515 136
rect -387 148 -384 151
rect -380 147 -377 150
rect -373 148 -370 151
rect -366 147 -363 150
rect -357 148 -354 151
rect -350 147 -347 150
rect -343 148 -340 151
rect -336 147 -333 150
rect -329 148 -326 151
rect -321 147 -318 150
rect -299 149 -296 152
rect -292 147 -289 150
rect -480 141 -477 144
rect -472 140 -469 143
rect -443 141 -440 144
rect -435 140 -432 143
rect -519 124 -515 128
rect -519 111 -515 115
rect -519 102 -515 106
rect -519 93 -515 97
rect -519 84 -515 88
rect -519 7 -515 11
rect -519 -1 -515 3
rect -519 -12 -515 -8
rect -404 4 -401 7
rect -397 3 -394 6
rect -390 4 -387 7
rect -383 3 -380 6
rect -374 4 -371 7
rect -367 3 -364 6
rect -360 4 -357 7
rect -353 3 -350 6
rect -346 4 -343 7
rect -338 3 -335 6
rect -316 5 -313 8
rect -309 3 -306 6
rect -480 -3 -477 0
rect -472 -4 -469 -1
rect -449 -3 -446 0
rect -441 -4 -438 -1
rect -519 -20 -515 -16
rect -519 -33 -515 -29
rect -519 -42 -515 -38
rect -519 -51 -515 -47
rect -519 -60 -515 -56
<< psubstratepcontact >>
rect -561 325 -557 329
rect -561 315 -557 319
rect -561 220 -557 224
rect -561 210 -557 214
rect -561 107 -557 111
rect -561 97 -557 101
rect -561 -37 -557 -33
rect -561 -47 -557 -43
<< nsubstratencontact >>
rect -506 325 -502 329
rect -506 315 -502 319
rect -506 220 -502 224
rect -506 210 -502 214
rect -506 107 -502 111
rect -506 97 -502 101
rect -506 -37 -502 -33
rect -506 -47 -502 -43
<< polysilicon >>
rect -554 378 -505 380
rect -554 368 -552 378
rect -571 366 -548 368
rect -542 366 -541 368
rect -539 366 -520 368
rect -513 366 -510 368
rect -571 295 -569 366
rect -539 349 -537 366
rect -507 349 -505 378
rect -476 362 -474 364
rect -476 352 -474 356
rect -566 347 -548 349
rect -542 347 -537 349
rect -524 347 -520 349
rect -513 347 -505 349
rect -500 349 -480 352
rect -475 349 -474 352
rect -476 348 -474 349
rect -566 309 -564 347
rect -476 343 -474 345
rect -534 327 -530 330
rect -555 325 -548 327
rect -542 325 -520 327
rect -513 325 -508 327
rect -533 317 -531 325
rect -534 309 -530 314
rect -566 307 -548 309
rect -542 307 -520 309
rect -513 307 -508 309
rect -571 293 -530 295
rect -510 286 -508 307
rect -472 307 -470 339
rect -342 332 -340 345
rect -435 328 -433 330
rect -393 328 -391 331
rect -375 328 -373 331
rect -435 318 -433 322
rect -393 319 -391 323
rect -434 315 -433 318
rect -425 316 -391 319
rect -435 314 -433 315
rect -393 312 -391 316
rect -375 315 -373 323
rect -342 322 -340 326
rect -341 319 -340 322
rect -342 318 -340 319
rect -381 313 -373 315
rect -342 313 -340 315
rect -381 312 -380 313
rect -375 312 -373 313
rect -435 309 -433 311
rect -393 308 -391 309
rect -472 305 -440 307
rect -381 286 -380 309
rect -375 308 -373 309
rect -510 284 -380 286
rect -554 273 -505 275
rect -554 263 -552 273
rect -571 261 -548 263
rect -542 261 -541 263
rect -539 261 -520 263
rect -513 261 -510 263
rect -571 190 -569 261
rect -539 244 -537 261
rect -507 244 -505 273
rect -476 257 -474 259
rect -476 247 -474 251
rect -566 242 -548 244
rect -542 242 -537 244
rect -524 242 -520 244
rect -513 242 -505 244
rect -500 244 -480 247
rect -475 244 -474 247
rect -476 243 -474 244
rect -566 204 -564 242
rect -350 242 -348 255
rect -476 238 -474 240
rect -437 238 -435 240
rect -401 238 -399 241
rect -383 238 -381 241
rect -534 222 -530 225
rect -555 220 -548 222
rect -542 220 -520 222
rect -513 220 -508 222
rect -533 212 -531 220
rect -476 217 -474 234
rect -309 238 -307 241
rect -437 228 -435 232
rect -401 229 -399 233
rect -436 225 -435 228
rect -425 226 -399 229
rect -437 224 -435 225
rect -401 222 -399 226
rect -383 225 -381 233
rect -350 232 -348 236
rect -349 229 -348 232
rect -339 230 -326 233
rect -350 228 -348 229
rect -329 229 -326 230
rect -309 229 -307 233
rect -389 223 -381 225
rect -329 226 -307 229
rect -350 223 -348 225
rect -389 222 -388 223
rect -383 222 -381 223
rect -309 222 -307 226
rect -299 225 -297 254
rect -258 242 -256 255
rect -291 238 -289 241
rect -211 237 -209 239
rect -205 237 -203 320
rect -201 237 -199 239
rect -191 237 -189 239
rect -181 237 -179 239
rect -167 237 -165 239
rect -291 225 -289 233
rect -258 232 -256 236
rect -257 229 -256 232
rect -258 228 -256 229
rect -211 229 -209 232
rect -299 223 -289 225
rect -205 229 -203 232
rect -201 229 -199 232
rect -191 230 -189 232
rect -205 227 -199 229
rect -258 223 -256 225
rect -291 222 -289 223
rect -211 222 -209 227
rect -201 222 -199 227
rect -191 222 -189 228
rect -181 230 -179 232
rect -181 222 -179 228
rect -167 227 -165 232
rect -166 225 -165 227
rect -167 222 -165 225
rect -437 219 -435 221
rect -401 218 -399 219
rect -476 215 -442 217
rect -534 204 -530 209
rect -389 204 -388 219
rect -383 218 -381 219
rect -309 218 -307 219
rect -291 218 -289 219
rect -211 218 -209 219
rect -201 218 -199 219
rect -191 218 -189 219
rect -181 218 -179 219
rect -167 218 -165 219
rect -566 202 -548 204
rect -542 202 -520 204
rect -513 202 -388 204
rect -571 188 -530 190
rect -554 160 -505 162
rect -554 150 -552 160
rect -571 148 -548 150
rect -542 148 -541 150
rect -539 148 -520 150
rect -513 148 -510 150
rect -571 77 -569 148
rect -539 131 -537 148
rect -507 131 -505 160
rect -383 152 -381 153
rect -369 152 -367 153
rect -353 152 -351 153
rect -339 152 -337 153
rect -324 152 -322 153
rect -295 152 -293 153
rect -476 144 -474 146
rect -439 144 -437 146
rect -383 140 -381 146
rect -476 134 -474 138
rect -439 134 -437 138
rect -382 137 -381 140
rect -369 138 -367 146
rect -353 138 -351 146
rect -339 138 -337 146
rect -324 138 -322 146
rect -295 142 -293 146
rect -566 129 -548 131
rect -542 129 -537 131
rect -524 129 -520 131
rect -513 129 -505 131
rect -500 131 -480 134
rect -475 131 -474 134
rect -438 131 -437 134
rect -383 132 -381 137
rect -369 132 -367 135
rect -353 132 -351 135
rect -339 132 -337 135
rect -324 132 -322 135
rect -295 132 -293 139
rect -476 130 -474 131
rect -439 130 -437 131
rect -566 91 -564 129
rect -476 125 -474 127
rect -383 128 -381 129
rect -369 128 -367 129
rect -353 128 -351 129
rect -339 128 -337 129
rect -324 128 -322 129
rect -295 128 -293 129
rect -439 125 -437 127
rect -470 121 -443 123
rect -439 121 -438 123
rect -534 109 -530 112
rect -555 107 -548 109
rect -542 107 -520 109
rect -513 107 -508 109
rect -528 100 -526 107
rect -534 95 -530 96
rect -534 92 -533 95
rect -531 92 -530 95
rect -534 91 -530 92
rect -566 89 -548 91
rect -542 89 -520 91
rect -513 89 -508 91
rect -571 75 -530 77
rect -554 16 -505 18
rect -554 6 -552 16
rect -571 4 -548 6
rect -542 4 -541 6
rect -539 4 -520 6
rect -513 4 -510 6
rect -571 -67 -569 4
rect -539 -13 -537 4
rect -507 -13 -505 16
rect -400 8 -398 9
rect -386 8 -384 9
rect -370 8 -368 9
rect -356 8 -354 9
rect -341 8 -339 9
rect -312 8 -310 9
rect -476 0 -474 2
rect -445 0 -443 2
rect -400 -4 -398 2
rect -476 -10 -474 -6
rect -445 -10 -443 -6
rect -399 -7 -398 -4
rect -386 -6 -384 2
rect -370 -6 -368 2
rect -356 -6 -354 2
rect -341 -6 -339 2
rect -312 -2 -310 2
rect -566 -15 -548 -13
rect -542 -15 -537 -13
rect -524 -15 -520 -13
rect -513 -15 -505 -13
rect -500 -13 -480 -10
rect -475 -13 -474 -10
rect -444 -13 -443 -10
rect -400 -12 -398 -7
rect -386 -12 -384 -9
rect -370 -12 -368 -9
rect -356 -12 -354 -9
rect -341 -12 -339 -9
rect -312 -12 -310 -5
rect -476 -14 -474 -13
rect -445 -14 -443 -13
rect -566 -53 -564 -15
rect -476 -19 -474 -17
rect -400 -16 -398 -15
rect -386 -16 -384 -15
rect -370 -16 -368 -15
rect -356 -16 -354 -15
rect -341 -16 -339 -15
rect -312 -16 -310 -15
rect -445 -19 -443 -17
rect -534 -35 -530 -32
rect -555 -37 -548 -35
rect -542 -37 -520 -35
rect -513 -37 -508 -35
rect -528 -43 -526 -37
rect -534 -49 -530 -48
rect -534 -51 -533 -49
rect -531 -51 -530 -49
rect -534 -53 -530 -51
rect -566 -55 -548 -53
rect -542 -55 -520 -53
rect -513 -55 -508 -53
rect -571 -69 -530 -67
<< polycontact >>
rect -503 348 -500 352
rect -480 349 -475 352
rect -473 339 -470 341
rect -534 330 -530 334
rect -533 315 -531 317
rect -534 295 -530 299
rect -437 315 -434 318
rect -428 316 -425 319
rect -344 319 -341 322
rect -206 320 -203 323
rect -440 305 -437 307
rect -503 243 -500 247
rect -480 244 -475 247
rect -299 254 -297 260
rect -476 234 -474 236
rect -534 225 -530 229
rect -439 225 -436 228
rect -430 226 -425 229
rect -352 229 -349 232
rect -343 230 -339 233
rect -260 229 -257 232
rect -211 227 -209 229
rect -192 228 -189 230
rect -181 228 -179 230
rect -167 225 -166 227
rect -442 215 -437 217
rect -533 210 -531 212
rect -534 190 -530 194
rect -385 137 -382 140
rect -296 139 -293 142
rect -503 130 -500 134
rect -480 131 -475 134
rect -441 131 -438 134
rect -370 135 -367 138
rect -354 135 -351 138
rect -340 135 -337 138
rect -325 135 -322 138
rect -474 121 -470 123
rect -443 121 -439 123
rect -534 112 -530 116
rect -528 98 -526 100
rect -533 92 -531 95
rect -534 77 -530 81
rect -402 -7 -399 -4
rect -313 -5 -310 -2
rect -503 -14 -500 -10
rect -480 -13 -475 -10
rect -447 -13 -444 -10
rect -387 -9 -384 -6
rect -371 -9 -368 -6
rect -357 -9 -354 -6
rect -342 -9 -339 -6
rect -534 -32 -530 -28
rect -528 -46 -526 -43
rect -533 -51 -531 -49
rect -534 -67 -530 -63
<< metal1 >>
rect -543 369 -519 373
rect -515 369 -495 373
rect -543 361 -519 365
rect -515 361 -500 365
rect -561 350 -547 354
rect -543 350 -519 354
rect -504 352 -500 361
rect -561 339 -557 350
rect -504 348 -503 352
rect -504 346 -500 348
rect -543 342 -519 346
rect -515 342 -500 346
rect -499 339 -495 369
rect -561 335 -536 339
rect -561 329 -547 333
rect -561 323 -557 325
rect -540 324 -536 335
rect -534 335 -495 339
rect -491 368 -459 370
rect -534 334 -530 335
rect -515 329 -502 333
rect -579 321 -557 323
rect -579 289 -577 321
rect -561 319 -557 321
rect -543 320 -519 324
rect -506 323 -502 325
rect -491 323 -488 368
rect -481 367 -477 368
rect -480 362 -477 367
rect -472 353 -469 358
rect -472 350 -465 353
rect -472 348 -469 350
rect -480 341 -477 344
rect -506 320 -488 323
rect -483 339 -473 341
rect -506 319 -502 320
rect -531 315 -528 317
rect -561 311 -547 315
rect -515 311 -502 315
rect -543 302 -519 306
rect -534 299 -530 302
rect -483 289 -481 339
rect -579 287 -481 289
rect -461 335 -459 368
rect -346 338 -335 339
rect -346 335 -343 338
rect -461 333 -343 335
rect -579 218 -577 287
rect -543 264 -519 268
rect -515 264 -495 268
rect -461 265 -459 333
rect -439 328 -436 333
rect -396 327 -394 333
rect -379 327 -377 333
rect -346 332 -343 333
rect -431 314 -428 324
rect -390 318 -388 324
rect -372 318 -370 325
rect -338 323 -335 328
rect -354 319 -344 322
rect -338 320 -206 323
rect -354 318 -352 319
rect -390 316 -352 318
rect -338 318 -335 320
rect -372 312 -370 316
rect -439 307 -436 310
rect -346 311 -343 314
rect -396 307 -394 309
rect -346 309 -335 311
rect -346 307 -342 309
rect -437 305 -342 307
rect -543 256 -519 260
rect -515 256 -500 260
rect -561 245 -547 249
rect -543 245 -519 249
rect -504 247 -500 256
rect -561 234 -557 245
rect -504 243 -503 247
rect -504 241 -500 243
rect -543 237 -519 241
rect -515 237 -500 241
rect -499 234 -495 264
rect -561 230 -536 234
rect -561 224 -547 228
rect -561 218 -557 220
rect -540 219 -536 230
rect -534 230 -495 234
rect -491 263 -459 265
rect -534 229 -530 230
rect -515 224 -502 228
rect -579 216 -557 218
rect -579 184 -577 216
rect -561 214 -557 216
rect -543 215 -519 219
rect -506 218 -502 220
rect -491 218 -488 263
rect -481 262 -477 263
rect -480 257 -477 262
rect -472 248 -469 253
rect -472 245 -466 248
rect -461 245 -459 263
rect -299 260 -297 270
rect -354 248 -343 249
rect -262 248 -213 250
rect -354 245 -351 248
rect -262 245 -259 248
rect -472 243 -469 245
rect -461 243 -259 245
rect -480 236 -477 239
rect -506 215 -488 218
rect -483 234 -476 236
rect -474 234 -470 236
rect -506 214 -502 215
rect -531 210 -528 212
rect -561 206 -547 210
rect -515 206 -502 210
rect -543 197 -519 201
rect -534 194 -530 197
rect -483 184 -481 234
rect -579 182 -481 184
rect -579 105 -577 182
rect -461 159 -459 243
rect -441 238 -438 243
rect -404 237 -402 243
rect -387 237 -385 243
rect -354 242 -351 243
rect -433 224 -430 234
rect -398 228 -396 234
rect -380 228 -378 235
rect -362 229 -352 232
rect -362 228 -360 229
rect -398 226 -360 228
rect -346 228 -343 238
rect -312 237 -310 243
rect -295 237 -293 243
rect -262 242 -259 243
rect -215 242 -213 248
rect -380 222 -378 226
rect -441 217 -438 220
rect -306 228 -304 234
rect -288 228 -286 235
rect -254 233 -251 238
rect -215 240 -165 242
rect -215 236 -213 240
rect -170 236 -168 240
rect -270 229 -260 232
rect -254 230 -231 233
rect -270 228 -268 229
rect -306 226 -268 228
rect -254 228 -251 230
rect -354 221 -351 224
rect -288 222 -286 226
rect -404 217 -402 219
rect -354 219 -343 221
rect -233 229 -231 230
rect -233 227 -211 229
rect -178 227 -176 233
rect -164 227 -162 233
rect -208 225 -167 227
rect -164 225 -159 227
rect -262 221 -259 224
rect -208 222 -206 225
rect -198 222 -196 225
rect -188 222 -186 225
rect -178 222 -176 225
rect -164 222 -162 225
rect -354 217 -350 219
rect -312 217 -310 219
rect -262 219 -251 221
rect -262 217 -258 219
rect -215 217 -213 220
rect -204 217 -202 220
rect -194 217 -192 220
rect -184 217 -182 220
rect -170 217 -168 220
rect -437 215 -168 217
rect -461 156 -295 159
rect -543 151 -519 155
rect -515 151 -495 155
rect -461 152 -459 156
rect -543 143 -519 147
rect -515 143 -500 147
rect -561 132 -547 136
rect -543 132 -519 136
rect -504 134 -500 143
rect -561 121 -557 132
rect -504 130 -503 134
rect -504 128 -500 130
rect -543 124 -519 128
rect -515 124 -500 128
rect -499 121 -495 151
rect -561 117 -536 121
rect -561 111 -547 115
rect -561 105 -557 107
rect -540 106 -536 117
rect -534 117 -495 121
rect -491 151 -459 152
rect -387 151 -384 156
rect -491 150 -432 151
rect -534 116 -530 117
rect -515 111 -502 115
rect -579 103 -557 105
rect -579 71 -577 103
rect -561 101 -557 103
rect -543 102 -519 106
rect -506 105 -502 107
rect -491 105 -488 150
rect -481 149 -477 150
rect -480 144 -477 149
rect -461 149 -440 150
rect -472 130 -469 140
rect -480 123 -477 126
rect -506 102 -488 105
rect -483 121 -474 123
rect -506 101 -502 102
rect -561 93 -547 97
rect -528 96 -526 98
rect -515 93 -502 97
rect -543 84 -519 88
rect -534 81 -530 84
rect -483 71 -481 121
rect -579 69 -481 71
rect -579 -39 -577 69
rect -461 15 -459 149
rect -443 144 -440 149
rect -373 151 -370 156
rect -357 151 -354 156
rect -380 142 -377 147
rect -343 151 -340 156
rect -366 142 -363 147
rect -329 151 -326 156
rect -350 142 -347 147
rect -299 152 -296 156
rect -336 142 -333 147
rect -321 142 -318 147
rect -292 142 -289 147
rect -195 142 -193 181
rect -435 135 -432 140
rect -410 137 -385 140
rect -380 139 -296 142
rect -292 139 -193 142
rect -410 135 -408 137
rect -343 135 -340 138
rect -435 132 -408 135
rect -318 132 -315 139
rect -292 132 -289 139
rect -435 130 -432 132
rect -443 123 -440 126
rect -387 124 -384 129
rect -299 124 -296 129
rect -387 123 -296 124
rect -444 121 -443 123
rect -439 121 -296 123
rect -461 12 -312 15
rect -543 7 -519 11
rect -515 7 -495 11
rect -461 8 -459 12
rect -543 -1 -519 3
rect -515 -1 -500 3
rect -561 -12 -547 -8
rect -543 -12 -519 -8
rect -504 -10 -500 -1
rect -561 -23 -557 -12
rect -504 -14 -503 -10
rect -504 -16 -500 -14
rect -543 -20 -519 -16
rect -515 -20 -500 -16
rect -499 -23 -495 7
rect -561 -27 -536 -23
rect -561 -33 -547 -29
rect -561 -39 -557 -37
rect -540 -38 -536 -27
rect -534 -27 -495 -23
rect -491 6 -438 8
rect -404 7 -401 12
rect -534 -28 -530 -27
rect -515 -33 -502 -29
rect -579 -41 -557 -39
rect -579 -73 -577 -41
rect -561 -43 -557 -41
rect -543 -42 -519 -38
rect -506 -39 -502 -37
rect -491 -39 -488 6
rect -481 5 -477 6
rect -450 5 -446 6
rect -480 0 -477 5
rect -449 0 -446 5
rect -390 7 -387 12
rect -374 7 -371 12
rect -472 -9 -469 -4
rect -397 -2 -394 3
rect -360 7 -357 12
rect -383 -2 -380 3
rect -346 7 -343 12
rect -367 -2 -364 3
rect -316 8 -313 12
rect -353 -2 -350 3
rect -338 -2 -335 3
rect -309 -2 -306 3
rect -185 -2 -183 135
rect -441 -9 -438 -4
rect -420 -7 -402 -4
rect -397 -5 -313 -2
rect -309 -5 -183 -2
rect -420 -9 -418 -7
rect -472 -12 -466 -9
rect -472 -14 -469 -12
rect -441 -12 -418 -9
rect -335 -12 -332 -5
rect -309 -12 -306 -5
rect -441 -14 -438 -12
rect -480 -21 -477 -18
rect -449 -21 -446 -18
rect -404 -20 -401 -15
rect -316 -20 -313 -15
rect -404 -21 -313 -20
rect -506 -42 -488 -39
rect -483 -23 -313 -21
rect -506 -43 -502 -42
rect -528 -47 -526 -46
rect -561 -51 -547 -47
rect -515 -51 -502 -47
rect -543 -60 -519 -56
rect -534 -63 -530 -60
rect -483 -73 -481 -23
rect -579 -75 -481 -73
<< m2contact >>
rect -528 315 -526 317
rect -440 315 -437 318
rect -528 210 -525 212
rect -441 225 -439 228
rect -195 228 -192 230
rect -183 228 -181 230
rect -195 181 -193 186
rect -528 92 -526 96
rect -533 90 -531 92
rect -373 135 -370 138
rect -443 131 -441 134
rect -185 135 -183 141
rect -450 -13 -447 -10
rect -528 -52 -526 -47
<< metal2 >>
rect -528 299 -526 315
rect -468 315 -440 318
rect -468 299 -466 315
rect -528 297 -466 299
rect -453 225 -441 228
rect -527 195 -525 210
rect -453 195 -451 225
rect -527 193 -451 195
rect -195 186 -193 228
rect -185 141 -183 230
rect -454 131 -443 134
rect -533 81 -531 90
rect -528 81 -526 92
rect -454 81 -452 131
rect -534 77 -530 81
rect -528 79 -452 81
rect -533 66 -531 77
rect -375 66 -373 138
rect -533 64 -373 66
rect -460 -13 -450 -10
rect -528 -63 -526 -52
rect -460 -63 -458 -13
rect -528 -65 -458 -63
<< m123contact >>
rect -465 350 -463 353
rect -299 270 -297 275
rect -466 245 -463 248
rect -469 132 -466 135
rect -357 135 -354 138
rect -328 135 -325 138
rect -390 -9 -387 -6
rect -374 -9 -371 -6
rect -360 -9 -357 -6
rect -345 -9 -342 -6
rect -533 -54 -531 -51
<< metal3 >>
rect -465 277 -463 350
rect -465 275 -297 277
rect -465 188 -463 245
rect -465 186 -359 188
rect -361 138 -359 186
rect -325 169 -323 275
rect -333 167 -323 169
rect -333 138 -331 167
rect -361 135 -357 138
rect -333 135 -328 138
rect -466 132 -462 135
rect -464 29 -462 132
rect -361 29 -359 135
rect -464 27 -394 29
rect -396 -6 -394 27
rect -380 27 -359 29
rect -380 -6 -378 27
rect -333 24 -331 135
rect -363 22 -331 24
rect -363 -6 -361 22
rect -396 -9 -390 -6
rect -380 -9 -374 -6
rect -363 -9 -360 -6
rect -350 -9 -345 -6
rect -533 -83 -531 -54
rect -350 -83 -348 -9
rect -533 -85 -348 -83
<< labels >>
rlabel metal1 -520 -74 -520 -74 1 gnd
rlabel metal1 -489 6 -489 6 1 vdd
rlabel metal1 -467 -10 -467 -10 1 x0
rlabel m123contact -468 134 -468 134 1 x1
rlabel metal1 -467 247 -467 247 1 x2
rlabel metal1 -468 352 -468 352 1 x3
rlabel metal1 -341 136 -341 136 1 temp
rlabel polysilicon -532 327 -532 327 1 a3
rlabel polysilicon -532 311 -532 311 1 b3
rlabel metal1 -429 317 -429 317 1 a3_not
rlabel metal1 -336 322 -336 322 1 AlessB_3
rlabel polysilicon -532 207 -532 207 1 b2
rlabel polysilicon -532 222 -532 222 1 a2
rlabel metal1 -431 228 -431 228 1 a2_not
rlabel metal1 -252 232 -252 232 1 AlessB_2
rlabel metal1 -162 226 -162 226 7 AlessB
rlabel polysilicon -532 110 -532 110 1 a1
rlabel polysilicon -536 90 -536 90 1 b1
rlabel metal1 -433 134 -433 134 1 a1_not
rlabel metal1 -290 140 -290 140 1 AlessB_1
rlabel polysilicon -533 -34 -533 -34 1 a0
rlabel polysilicon -536 -54 -536 -54 1 b0
rlabel metal1 -438 -10 -438 -10 1 a0_not
rlabel metal1 -306 -4 -306 -4 1 AlessB_0
<< end >>
