* SPICE3 file created from final_1.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param width_P=8*LAMBDA
.param  width_N = 4*LAMBDA
.global gnd vdd
* .option scale=0.81u

Vdd vdd gnd 'SUPPLY'

* Vs0 s0 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
* Vs1 s1 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)

* Vs0 s0 gnd DC 1.8
* Vs1 s1 gnd DC 1.8

Vd0 D0 gnd DC 1.8
Vd1 D1 gnd DC 0
Vd2 D2 gnd DC 0
Vd3 D3 gnd DC 0

Va3 a3 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
Va2 a2 gnd PULSE(1.8 0 100ns 100ps 100ps 100ns 200ns)
Va1 a1 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
Va0 a0 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)

Vb3 b3 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
Vb2 b2 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)
Vb1 b1 gnd PULSE(1.8 0 200ns 100ps 100ps 200ns 400ns)
Vb0 b0 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)

.option scale=0.01u

M1000 D1 a_290_124# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=6.77095e+06 ps=89262
M1001 a_386_n38# D3 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1002 a_413_308# D0 a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1944 as=0 ps=0
M1003 a_476_230# a_437_308# a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1004 a_386_n184# a0 a_386_n198# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1005 a_381_n331# b2 a_246_106# w_371_n334# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=1.64353e+07 ps=162162
M1006 a_696_n179# b0 a_696_n193# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1007 comp_b1 a_696_n120# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1008 a_696_n120# b1 a_246_106# w_686_n123# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1009 a_476_574# b1 a_246_106# w_466_571# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1010 a_571_n426# and_b0 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1011 and_b1 a_381_n377# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1012 a_696_n179# D2 a_246_106# w_686_n182# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1013 a_476_404# a3 a_476_390# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1014 and_a2 a_386_n79# a_246_106# w_428_n78# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1015 D1 a_290_124# a_246_106# w_332_125# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1016 a_571_n316# and_b2 a_246_106# w_561_n319# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1017 a_476_244# a_491_234# a_246_106# w_466_241# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1018 and_a1 a_386_n125# a_246_106# w_428_n124# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1019 a_381_n276# b3 a_381_n290# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1020 a_696_n74# b2 a_696_n88# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1021 comp_a0 a_565_17# a_246_106# w_607_18# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1022 a_565_17# D2 a_246_106# w_555_14# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1023 and_oper_out1 a_571_n360# a_246_106# w_613_n359# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1024 a_386_n139# D3 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1025 a_476_574# a_437_308# a_246_106# w_466_571# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1026 a_290_75# s0_not a_246_106# w_280_72# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1027 and_a3 a_386_n24# a_246_106# w_428_n23# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1028 a_696_n134# D2 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1029 a_476_390# a_437_308# a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1030 a_386_n79# D3 a_246_106# w_376_n82# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1031 a_381_n450# D3 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1032 adsub_b1 a_476_574# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1033 a_571_n374# and_b1 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1034 a_571_n412# and_a0 a_571_n426# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1035 a_696_n19# b3 a_696_n33# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1036 a_476_244# a_437_308# a_246_106# w_466_241# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1037 adsub_a0 a_476_244# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1038 a_571_n316# and_a2 a_246_106# w_561_n319# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1039 a_381_n276# D3 a_246_106# w_371_n279# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1040 adsub_b1 a_476_574# a_246_106# w_518_575# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1041 a_386_n24# D3 a_246_106# w_376_n27# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1042 and_oper_out3 a_571_n263# a_246_106# w_613_n262# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1043 a_565_17# a0 a_246_106# w_555_14# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1044 a_413_321# D0 a_246_106# w_404_319# CMOSP w=405 l=162
+  ad=262440 pd=2106 as=0 ps=0
M1045 and_a0 a_386_n184# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1046 a_386_n184# a0 a_246_106# w_376_n187# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1047 a_476_404# a3 a_246_106# w_466_401# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1048 adsub_a0 a_476_244# a_246_106# w_518_245# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1049 a_381_n436# b0 a_381_n450# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1050 a_571_n412# and_b0 a_246_106# w_561_n415# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1051 a_571_n360# and_a1 a_571_n374# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1052 and_oper_out2 a_571_n316# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1053 a_571_n277# and_b3 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1054 comp_b2 a_696_n74# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1055 a_565_17# a0 a_565_3# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1056 adsub_a3 a_476_404# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1057 a_290_15# s1 a_246_95# Gnd CMOSN w=243 l=162
+  ad=216513 pd=2268 as=0 ps=0
M1058 a_696_n74# b2 a_246_106# w_686_n77# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1059 a_381_n276# b3 a_246_106# w_371_n279# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1060 D2 a_290_75# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1061 a_476_404# a_437_308# a_246_106# w_466_401# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1062 a_386_n125# D3 a_246_106# w_376_n128# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1063 comp_b1 a_696_n120# a_246_106# w_738_n119# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1064 a_290_176# s1_not a_290_162# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1065 and_b1 a_381_n377# a_246_106# w_423_n376# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1066 a_386_n79# a2 a_386_n93# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1067 a_381_n436# D3 a_246_106# w_371_n439# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1068 s0_not s0 a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1069 a_476_349# a2 a_476_335# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1070 s1_not s1 a_246_106# w_244_81# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1071 and_b2 a_381_n331# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1072 adsub_a2 a_476_349# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1073 D2 a_290_75# a_246_106# w_332_76# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1074 a_571_n412# and_a0 a_246_106# w_561_n415# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1075 a_290_75# s1 a_305_61# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=19683 ps=648
M1076 D3 a_290_29# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1077 a_571_n263# and_a3 a_571_n277# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1078 and_b3 a_381_n276# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1079 a_437_308# a_413_308# a_246_95# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1080 a_381_n391# D3 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1081 adsub_a3 a_476_404# a_246_106# w_518_405# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1082 a_565_62# D2 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1083 a_696_n88# D2 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1084 adsub_a2 a_476_349# a_246_106# w_518_350# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1085 a_565_177# a3 a_565_163# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1086 D3 a_290_29# a_246_106# w_332_30# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1087 a_476_515# b0 a_476_501# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1088 a_476_335# a_437_308# a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1089 a_290_29# s1 a_246_106# w_280_26# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1090 a_381_n436# b0 a_246_106# w_371_n439# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1091 a_571_n263# and_b3 a_246_106# w_561_n266# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1092 a_290_176# s1_not a_246_106# w_280_173# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1093 comp_b0 a_696_n179# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1094 a_696_n179# b0 a_246_106# w_686_n182# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1095 a_290_124# s1_not a_290_110# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1096 comp_a3 a_565_177# a_246_106# w_607_178# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1097 a_381_n377# b1 a_381_n391# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1098 a_696_n33# D2 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1099 a_476_349# a2 a_246_106# w_466_346# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1100 a_565_163# D2 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1101 a_290_75# s1 a_246_106# w_280_72# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1102 and_a0 a_386_n184# a_246_106# w_428_n183# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1103 a_476_501# a_437_308# a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1104 a_565_76# a1 a_565_62# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1105 a_565_76# D2 a_246_106# w_555_73# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1106 s1_not s1 a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1107 and_b0 a_381_n436# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1108 a_476_675# b3 a_476_661# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1109 and_oper_out2 a_571_n316# a_246_106# w_613_n315# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1110 comp_b2 a_696_n74# a_246_106# w_738_n73# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1111 a_386_n198# D3 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1112 a_386_n125# a1 a_386_n139# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1113 a_476_303# a1 a_246_106# w_466_300# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1114 a_565_177# a3 a_246_106# w_555_174# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1115 a_696_n193# D2 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1116 a_696_n120# b1 a_696_n134# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1117 a_696_n120# D2 a_246_106# w_686_n123# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1118 comp_b3 a_696_n19# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1119 a_476_515# b0 a_246_106# w_466_512# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1120 a_571_n263# and_a3 a_246_106# w_561_n266# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1121 a_476_349# a_437_308# a_246_106# w_466_346# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1122 a_437_308# a_413_308# a_246_106# w_404_319# CMOSP w=405 l=162
+  ad=131220 pd=1458 as=0 ps=0
M1123 a_571_n360# and_b1 a_246_106# w_561_n363# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1124 a_696_n19# b3 a_246_106# w_686_n22# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1125 a_476_303# a1 a_476_289# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1126 adsub_a1 a_476_303# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1127 a_696_n74# D2 a_246_106# w_686_n77# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1128 a_476_661# a_437_308# a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1129 a_290_124# s1_not a_246_106# w_280_121# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1130 and_b2 a_381_n331# a_246_106# w_423_n330# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1131 a_565_122# a2 a_246_106# w_555_119# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1132 a_386_n24# a3 a_386_n38# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1133 a_476_303# a_437_308# a_246_106# w_466_300# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1134 a_565_177# D2 a_246_106# w_555_174# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1135 a_476_515# a_437_308# a_246_106# w_466_512# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1136 comp_a3 a_565_177# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1137 s0_not s0 a_246_106# w_243_117# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1138 a_565_76# a1 a_246_106# w_555_73# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1139 and_oper_out3 a_571_n263# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1140 a_386_n93# D3 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1141 a_290_162# s0_not a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1142 and_b3 a_381_n276# a_246_106# w_423_n275# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1143 adsub_b0 a_476_515# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1144 a_290_29# s0 a_303_15# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=59049 ps=972
M1145 a_476_675# b3 a_246_106# w_466_672# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1146 and_oper_out0 a_571_n412# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1147 a_381_n345# D3 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1148 a_476_289# a_437_308# a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1149 a_571_n360# and_a1 a_246_106# w_561_n363# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1150 a_413_308# D1 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1151 comp_a1 a_565_76# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1152 adsub_a1 a_476_303# a_246_106# w_518_304# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1153 a_565_122# D2 a_246_106# w_555_119# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1154 adsub_b0 a_476_515# a_246_106# w_518_516# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1155 comp_a2 a_565_122# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1156 a_565_122# a2 a_565_108# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1157 and_a2 a_386_n79# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1158 a_476_620# b2 a_246_106# w_466_617# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1159 and_a1 a_386_n125# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1160 a_386_n125# a1 a_246_106# w_376_n128# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1161 comp_a1 a_565_76# a_246_106# w_607_77# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1162 comp_b0 a_696_n179# a_246_106# w_738_n178# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1163 a_386_n184# D3 a_246_106# w_376_n187# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1164 a_476_675# a_437_308# a_246_106# w_466_672# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1165 a_386_n79# a2 a_246_106# w_376_n82# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1166 adsub_b3 a_476_675# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1167 a_303_15# s0 a_290_15# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1168 and_oper_out1 a_571_n360# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1169 comp_a0 a_565_17# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1170 comp_a2 a_565_122# a_246_106# w_607_123# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1171 a_381_n331# b2 a_381_n345# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1172 a_290_176# s0_not a_246_106# w_280_173# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1173 and_a3 a_386_n24# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1174 D0 a_290_176# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1175 a_290_110# s0 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1176 a_565_108# D2 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1177 a_290_29# s0 a_246_106# w_280_26# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1178 a_565_3# D2 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1179 a_305_61# s1 a_290_61# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=255879 ps=2592
M1180 and_b0 a_381_n436# a_246_106# w_423_n435# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1181 a_381_n377# D3 a_246_106# w_371_n380# CMOSP w=405 l=162
+  ad=360855 pd=3402 as=0 ps=0
M1182 a_571_n330# and_b2 a_246_95# Gnd CMOSN w=243 l=162
+  ad=314928 pd=3078 as=0 ps=0
M1183 adsub_b3 a_476_675# a_246_106# w_518_676# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1184 a_476_620# a_437_308# a_246_106# w_466_617# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1185 a_386_n24# a3 a_246_106# w_376_n27# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1186 comp_b3 a_696_n19# a_246_106# w_738_n18# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1187 adsub_b2 a_476_620# a_246_95# Gnd CMOSN w=243 l=162
+  ad=118098 pd=1458 as=0 ps=0
M1188 a_476_620# b2 a_476_606# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1189 a_476_574# b1 a_476_560# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=314928 ps=3078
M1190 D0 a_290_176# a_246_106# w_332_177# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1191 a_381_n331# D3 a_246_106# w_371_n334# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1192 a_413_308# D1 a_413_321# w_404_319# CMOSP w=405 l=162
+  ad=98415 pd=1296 as=0 ps=0
M1193 a_476_244# a_491_234# a_476_230# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1194 adsub_b2 a_476_620# a_246_106# w_518_621# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
M1195 a_381_n377# b1 a_246_106# w_371_n380# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1196 a_696_n19# D2 a_246_106# w_686_n22# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1197 a_476_606# a_437_308# a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1198 a_571_n316# and_a2 a_571_n330# Gnd CMOSN w=243 l=162
+  ad=78732 pd=1134 as=0 ps=0
M1199 a_381_n290# D3 a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1200 a_290_124# s0 a_246_106# w_280_121# CMOSP w=405 l=162
+  ad=0 pd=0 as=0 ps=0
M1201 a_476_560# a_437_308# a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1202 a_290_61# s0_not a_246_95# Gnd CMOSN w=243 l=162
+  ad=0 pd=0 as=0 ps=0
M1203 and_oper_out0 a_571_n412# a_246_106# w_613_n411# CMOSP w=486 l=162
+  ad=236196 pd=1944 as=0 ps=0
C0 D1 a1 0.04fF
C1 w_686_n77# a_696_n74# 0.42fF
C2 w_518_245# a_246_106# 1.86fF
C3 a_476_574# b1 0.60fF
C4 a_246_106# a_386_n24# 0.60fF
C5 a1 D2 0.08fF
C6 w_555_119# a_246_106# 0.28fF
C7 w_466_241# a_437_308# 0.93fF
C8 w_738_n178# comp_b0 0.19fF
C9 w_466_401# a_246_106# 0.28fF
C10 w_561_n266# a_571_n263# 0.42fF
C11 w_428_n78# and_a2 0.19fF
C12 w_466_346# a_437_308# 0.93fF
C13 w_686_n77# D2 0.93fF
C14 w_376_n128# a1 1.08fF
C15 D2 a0 0.07fF
C16 w_607_178# comp_a3 0.19fF
C17 a_476_404# a_246_106# 0.60fF
C18 w_466_241# a_476_244# 0.42fF
C19 s1_not a_290_110# 0.06fF
C20 b3 a_696_n19# 0.87fF
C21 a0 a_565_17# 0.60fF
C22 a2 a_246_95# 1.38fF
C23 D0 a_246_106# 1.04fF
C24 w_555_73# a1 0.93fF
C25 w_518_304# adsub_a1 0.19fF
C26 w_738_n18# comp_b3 0.19fF
C27 a_246_95# a_491_234# 0.64fF
C28 s0_not a_246_95# 0.46fF
C29 w_243_117# a_246_106# 0.89fF
C30 a1 a_476_289# 0.06fF
C31 w_561_n415# and_b0 0.93fF
C32 b3 D2 0.64fF
C33 a1 a_246_95# 1.62fF
C34 w_466_617# a_246_106# 0.28fF
C35 w_607_18# a_565_17# 2.17fF
C36 w_613_n315# a_246_106# 1.14fF
C37 w_686_n22# b2 0.47fF
C38 a_476_675# b3 0.80fF
C39 w_371_n439# a_246_106# 0.28fF
C40 a_246_106# a_571_n263# 0.41fF
C41 w_371_n334# b2 2.12fF
C42 w_466_300# a1 0.93fF
C43 w_561_n415# and_a0 1.88fF
C44 w_466_672# b3 1.03fF
C45 and_a0 a_571_n412# 1.08fF
C46 w_376_n187# a_246_106# 0.28fF
C47 w_404_319# a_246_106# 2.54fF
C48 w_738_n119# a_246_106# 1.86fF
C49 a_246_95# a0 1.70fF
C50 a1 a_386_n139# 0.06fF
C51 w_428_n183# and_a0 0.19fF
C52 w_332_76# a_246_106# 1.79fF
C53 w_555_174# a3 1.09fF
C54 w_371_n279# a_246_106# 0.28fF
C55 and_a1 and_b3 0.27fF
C56 w_428_n23# a_246_106# 1.86fF
C57 w_555_174# D2 0.93fF
C58 b3 a_246_95# 2.10fF
C59 a_246_95# and_a1 0.27fF
C60 w_371_n439# b0 0.93fF
C61 a_246_106# a_476_574# 0.60fF
C62 b3 b1 0.27fF
C63 s0_not s1_not 4.30fF
C64 b3 and_a0 0.07fF
C65 and_a1 and_a0 0.82fF
C66 and_a2 and_b3 0.60fF
C67 w_518_676# adsub_b3 0.19fF
C68 w_423_n330# a_381_n331# 2.17fF
C69 w_423_n435# a_381_n436# 2.17fF
C70 w_280_121# a_290_124# 0.42fF
C71 w_686_n182# a_246_106# 0.28fF
C72 w_738_n119# comp_b1 0.19fF
C73 w_466_401# a_437_308# 0.93fF
C74 a_246_95# and_a2 0.46fF
C75 and_a2 and_a0 0.13fF
C76 a_246_106# a_565_177# 0.60fF
C77 w_686_n182# a_696_n179# 0.42fF
C78 w_518_245# a_476_244# 2.17fF
C79 b2 D3 0.07fF
C80 a_246_95# and_a3 0.60fF
C81 w_423_n275# a_381_n276# 2.17fF
C82 a2 a_246_106# 3.68fF
C83 a_246_106# a_381_n436# 0.60fF
C84 s0_not a_246_106# 0.73fF
C85 w_466_617# a_437_308# 0.93fF
C86 w_466_571# b1 0.93fF
C87 a1 a_246_106# 0.82fF
C88 w_686_n182# b0 0.93fF
C89 w_561_n415# a_246_106# 0.28fF
C90 a_246_106# a_381_n276# 0.60fF
C91 w_518_621# adsub_b2 0.19fF
C92 w_466_617# b2 2.12fF
C93 w_371_n380# b1 0.93fF
C94 w_466_512# a_246_106# 0.28fF
C95 a_246_106# a_571_n412# 0.41fF
C96 w_555_14# a0 0.93fF
C97 and_a1 and_b2 0.04fF
C98 w_428_n183# a_246_106# 2.31fF
C99 w_404_319# a_437_308# 0.14fF
C100 w_686_n77# a_246_106# 0.28fF
C101 a_246_106# a0 1.40fF
C102 w_428_n124# and_a1 0.19fF
C103 w_613_n262# and_oper_out3 0.19fF
C104 b2 a_696_n88# 0.10fF
C105 w_607_77# a_565_76# 2.17fF
C106 w_613_n262# a_246_106# 1.14fF
C107 w_280_72# s0_not 0.93fF
C108 w_244_81# s1_not 0.19fF
C109 w_607_18# a_246_106# 1.86fF
C110 b0 a_381_n436# 0.60fF
C111 w_555_73# a_565_76# 0.42fF
C112 b1 a_696_n134# 0.06fF
C113 w_371_n334# D3 0.93fF
C114 a_476_349# a2 1.06fF
C115 b3 a_246_106# 1.61fF
C116 w_561_n266# and_a3 2.64fF
C117 a_246_106# and_a1 1.16fF
C118 w_376_n27# a3 1.09fF
C119 a3 D2 0.10fF
C120 w_466_512# b0 0.93fF
C121 a_246_106# a_571_n360# 0.41fF
C122 w_518_516# adsub_b0 0.19fF
C123 w_376_n82# a_246_106# 0.28fF
C124 w_280_173# s1_not 0.93fF
C125 s1_not a_290_124# 0.60fF
C126 w_243_117# s0 0.66fF
C127 b1 a_696_n120# 0.60fF
C128 a_476_303# a1 0.60fF
C129 w_423_n376# and_b1 0.19fF
C130 a_246_106# and_a2 2.41fF
C131 w_332_177# a_246_106# 1.79fF
C132 w_332_30# D3 0.19fF
C133 w_613_n411# a_571_n412# 2.17fF
C134 w_404_319# a_413_308# 0.96fF
C135 w_244_81# a_246_106# 1.83fF
C136 w_376_n187# a_386_n184# 0.42fF
C137 a_476_675# w_466_672# 0.42fF
C138 w_561_n319# and_b2 0.93fF
C139 w_555_174# a_246_106# 0.28fF
C140 a_246_106# and_a3 1.40fF
C141 a_476_515# a_246_106# 0.60fF
C142 b0 b3 0.41fF
C143 a3 a_246_95# 1.08fF
C144 a_246_106# a_381_n331# 0.60fF
C145 D1 a_246_95# 2.01fF
C146 w_466_571# a_246_106# 0.28fF
C147 w_613_n359# and_oper_out1 0.19fF
C148 w_555_73# D2 0.93fF
C149 w_607_123# a_565_122# 2.17fF
C150 w_518_575# a_476_574# 2.17fF
C151 a1 a_437_308# 0.04fF
C152 a_290_124# a_246_106# 0.60fF
C153 w_280_173# a_246_106# 0.28fF
C154 a_491_234# a_476_230# 0.10fF
C155 w_371_n380# a_246_106# 0.28fF
C156 w_518_621# a_476_620# 2.17fF
C157 a_246_95# D2 5.64fF
C158 w_561_n319# a_246_106# 0.28fF
C159 w_613_n315# a_571_n316# 2.17fF
C160 b1 D2 0.04fF
C161 w_466_512# a_437_308# 0.93fF
C162 w_466_401# a_476_404# 0.42fF
C163 w_466_241# a_491_234# 0.93fF
C164 w_613_n359# a_571_n360# 2.17fF
C165 w_332_177# a_290_176# 2.17fF
C166 a_476_244# a_491_234# 0.60fF
C167 w_466_346# a2 2.12fF
C168 w_244_81# s1 0.66fF
C169 w_518_350# adsub_a2 0.19fF
C170 w_423_n376# a_246_106# 1.86fF
C171 b2 a0 0.67fF
C172 w_686_n77# b2 2.12fF
C173 a_476_515# b0 0.60fF
C174 w_607_18# comp_a0 0.19fF
C175 w_607_178# a_565_177# 2.17fF
C176 w_280_26# a_246_106# 0.28fF
C177 w_371_n439# D3 0.93fF
C178 and_a0 and_b3 0.46fF
C179 w_332_125# a_290_124# 2.17fF
C180 a_246_106# a_565_76# 0.60fF
C181 w_280_26# a_290_29# 0.42fF
C182 b3 b2 0.41fF
C183 a_246_106# a_476_620# 0.60fF
C184 b2 and_a1 0.06fF
C185 w_428_n23# a_386_n24# 2.17fF
C186 a_246_95# b1 1.62fF
C187 w_518_516# a_476_515# 2.17fF
C188 w_428_n78# a_246_106# 1.86fF
C189 a_246_95# and_a0 0.46fF
C190 a_246_106# a_696_n120# 0.60fF
C191 s0_not s0 0.07fF
C192 w_280_173# a_290_176# 0.42fF
C193 s1_not a_290_162# 0.06fF
C194 w_280_121# s1_not 0.93fF
C195 b0 a_696_n193# 0.10fF
C196 w_376_n187# D3 0.93fF
C197 a0 a_386_n198# 0.10fF
C198 a_246_106# a_290_75# 0.60fF
C199 w_371_n279# D3 0.93fF
C200 b2 and_a2 0.46fF
C201 a_246_106# a_696_n74# 0.60fF
C202 w_518_350# a_246_106# 1.86fF
C203 w_404_319# D0 0.80fF
C204 w_428_n183# a_386_n184# 2.17fF
C205 a1 a_386_n125# 0.87fF
C206 a_386_n184# a0 1.06fF
C207 w_423_n330# and_b2 0.19fF
C208 a_246_106# a_565_122# 0.60fF
C209 w_280_26# s1 0.93fF
C210 a2 a_386_n79# 1.06fF
C211 b2 and_a3 0.60fF
C212 and_a0 and_b1 0.07fF
C213 a3 a_246_106# 1.89fF
C214 w_561_n266# and_b3 0.93fF
C215 a_246_106# a_696_n19# 0.60fF
C216 w_466_571# a_437_308# 0.93fF
C217 D1 a_246_106# 1.04fF
C218 w_555_14# D2 0.93fF
C219 w_280_72# a_290_75# 0.42fF
C220 b2 a_381_n331# 1.06fF
C221 s1_not a_246_95# 1.35fF
C222 w_280_121# a_246_106# 0.28fF
C223 w_376_n27# a_246_106# 0.28fF
C224 w_686_n22# b3 1.09fF
C225 w_423_n435# and_b0 0.19fF
C226 w_561_n363# and_a1 1.08fF
C227 a_246_106# D2 1.83fF
C228 w_555_14# a_565_17# 0.42fF
C229 w_423_n330# a_246_106# 1.86fF
C230 a_476_675# a_246_106# 0.60fF
C231 w_555_119# a2 2.12fF
C232 a_290_75# s1 0.60fF
C233 a_246_106# a_565_17# 0.60fF
C234 w_561_n363# a_571_n360# 0.42fF
C235 w_466_672# a_246_106# 0.28fF
C236 a_476_675# w_518_676# 2.17fF
C237 w_423_n275# and_b3 0.19fF
C238 w_518_350# a_476_349# 2.17fF
C239 w_518_304# a_246_106# 1.86fF
C240 w_376_n128# a_246_106# 0.28fF
C241 and_a0 and_b2 0.07fF
C242 w_686_n123# a_696_n120# 0.42fF
C243 w_607_77# a_246_106# 1.86fF
C244 a_246_106# and_b3 1.21fF
C245 a1 D3 0.04fF
C246 w_332_125# D1 0.19fF
C247 w_555_73# a_246_106# 0.28fF
C248 a_246_106# a_246_95# 0.87fF
C249 w_376_n82# a_386_n79# 0.42fF
C250 a_476_620# b2 1.06fF
C251 a_246_106# and_a0 1.47fF
C252 D0 a1 0.06fF
C253 w_466_300# a_246_106# 0.28fF
C254 w_243_117# s0_not 0.19fF
C255 w_371_n334# a_381_n331# 0.42fF
C256 w_371_n439# a_381_n436# 0.42fF
C257 w_607_77# comp_a1 0.19fF
C258 D3 a0 0.07fF
C259 w_607_123# a_246_106# 1.86fF
C260 w_518_405# a_246_106# 1.86fF
C261 a2 a_565_108# 0.10fF
C262 w_371_n380# a_381_n377# 0.42fF
C263 and_a2 a_571_n316# 1.21fF
C264 D0 a0 0.09fF
C265 b2 a_696_n74# 1.06fF
C266 b3 D3 0.06fF
C267 w_686_n123# D2 0.93fF
C268 a_246_106# and_b1 1.40fF
C269 w_738_n73# a_696_n74# 2.17fF
C270 w_518_304# a_476_303# 2.17fF
C271 w_423_n376# a_381_n377# 2.17fF
C272 w_376_n82# D3 0.93fF
C273 b0 a_246_95# 1.79fF
C274 a_246_95# s1 2.01fF
C275 w_613_n262# a_571_n263# 2.17fF
C276 w_371_n279# a_381_n276# 0.42fF
C277 b0 b1 1.23fF
C278 w_280_26# s0 0.93fF
C279 b2 a_696_n19# 0.46fF
C280 s1_not a_246_106# 0.27fF
C281 w_518_621# a_246_106# 1.86fF
C282 w_376_n187# a0 1.88fF
C283 w_561_n266# a_246_106# 0.28fF
C284 w_423_n435# a_246_106# 1.86fF
C285 b2 D2 0.07fF
C286 w_561_n319# a_571_n316# 0.42fF
C287 w_466_300# a_476_303# 0.42fF
C288 w_466_672# a_437_308# 0.93fF
C289 w_332_177# D0 0.19fF
C290 a_246_106# and_b2 1.40fF
C291 w_738_n178# a_246_106# 1.86fF
C292 w_428_n124# a_246_106# 1.86fF
C293 a2 a_565_177# 0.46fF
C294 w_607_123# comp_a2 0.19fF
C295 w_686_n123# b1 0.93fF
C296 w_423_n275# a_246_106# 1.86fF
C297 w_371_n279# b3 1.09fF
C298 b0 a_476_501# 0.10fF
C299 w_613_n315# and_oper_out2 0.19fF
C300 b2 and_b3 0.60fF
C301 w_518_575# adsub_b1 0.19fF
C302 w_371_n380# D3 0.93fF
C303 w_555_14# a_246_106# 0.28fF
C304 w_738_n178# a_696_n179# 2.17fF
C305 a1 a_565_62# 0.06fF
C306 a_437_308# a_246_95# 4.88fF
C307 b3 a_696_n33# 0.06fF
C308 w_428_n78# a_386_n79# 2.17fF
C309 D1 a_413_308# 0.60fF
C310 and_a3 a_571_n263# 1.21fF
C311 a0 a_565_3# 0.10fF
C312 a_246_95# b2 3.51fF
C313 a_437_308# b1 0.04fF
C314 w_686_n22# a_696_n19# 0.42fF
C315 a_290_176# s1_not 0.60fF
C316 a_246_106# a_290_29# 0.60fF
C317 w_466_300# a_437_308# 0.93fF
C318 b2 b1 0.46fF
C319 w_518_676# a_246_106# 1.86fF
C320 b2 and_a0 0.07fF
C321 w_280_121# s0 1.12fF
C322 a_246_106# a_696_n179# 0.60fF
C323 w_686_n22# D2 0.93fF
C324 w_738_n18# a_696_n19# 2.17fF
C325 w_561_n415# a_571_n412# 0.42fF
C326 w_280_72# a_246_106# 0.28fF
C327 w_428_n23# and_a3 0.19fF
C328 a1 a0 0.41fF
C329 w_332_125# a_246_106# 1.79fF
C330 a_476_349# a_246_106# 0.60fF
C331 a_476_560# b1 0.06fF
C332 b1 a_381_n391# 0.06fF
C333 a_290_176# a_246_106# 0.60fF
C334 w_555_119# a_565_122# 0.42fF
C335 w_376_n128# a_386_n125# 0.42fF
C336 w_466_571# a_476_574# 0.42fF
C337 a1 b3 0.31fF
C338 a_476_303# a_246_106# 0.60fF
C339 s0 a_246_95# 1.21fF
C340 w_376_n82# a2 2.12fF
C341 b0 a_696_n179# 0.60fF
C342 a3 a_386_n24# 0.87fF
C343 w_613_n411# a_246_106# 1.14fF
C344 b3 a_381_n276# 0.87fF
C345 w_466_617# a_476_620# 0.42fF
C346 w_613_n359# a_246_106# 1.14fF
C347 w_518_516# a_246_106# 1.86fF
C348 w_518_405# adsub_a3 0.19fF
C349 w_466_401# a3 1.09fF
C350 b1 a_381_n377# 0.60fF
C351 w_376_n27# a_386_n24# 0.42fF
C352 w_555_174# a_565_177# 0.42fF
C353 w_555_119# D2 0.93fF
C354 w_686_n123# a_246_106# 0.28fF
C355 a1 and_a2 0.41fF
C356 w_280_72# s1 0.93fF
C357 b3 a0 1.06fF
C358 and_a1 a0 0.27fF
C359 w_518_245# adsub_a0 0.19fF
C360 w_555_174# a2 0.47fF
C361 a2 and_a3 0.07fF
C362 w_738_n119# a_696_n120# 2.17fF
C363 a_476_404# a3 0.87fF
C364 w_376_n27# D3 0.93fF
C365 w_561_n363# and_b1 0.93fF
C366 a_437_308# a_246_106# 0.60fF
C367 a1 and_a3 0.04fF
C368 b3 and_a1 0.06fF
C369 and_a2 a0 0.46fF
C370 a_246_106# b2 3.51fF
C371 w_332_76# a_290_75# 2.17fF
C372 w_466_512# a_476_515# 0.42fF
C373 w_738_n73# a_246_106# 1.86fF
C374 s1_not s0 0.04fF
C375 w_280_173# s0_not 0.93fF
C376 and_a1 a_571_n360# 0.89fF
C377 w_376_n128# D3 0.93fF
C378 b3 and_a2 0.09fF
C379 w_466_241# a_246_106# 0.28fF
C380 and_a3 a0 0.07fF
C381 and_a2 and_a1 0.58fF
C382 a_246_106# a_476_244# 0.60fF
C383 w_466_346# a_246_106# 0.28fF
C384 w_404_319# D1 0.80fF
C385 a_246_95# D3 5.44fF
C386 b1 D3 0.04fF
C387 b3 and_a3 0.60fF
C388 and_a3 and_a1 0.10fF
C389 b0 a_437_308# 0.07fF
C390 w_332_76# D2 0.19fF
C391 b0 b2 0.46fF
C392 b0 a_381_n450# 0.10fF
C393 w_518_575# a_246_106# 1.86fF
C394 a_246_106# a_386_n184# 0.60fF
C395 w_428_n124# a_386_n125# 2.17fF
C396 w_607_178# a_246_106# 1.86fF
C397 s0 a_246_106# 0.60fF
C398 a1 a_565_76# 0.60fF
C399 w_686_n22# a_246_106# 0.28fF
C400 w_561_n363# a_246_106# 0.28fF
C401 a3 a_565_163# 0.06fF
C402 and_a3 and_a2 0.16fF
C403 w_371_n334# a_246_106# 0.28fF
C404 a_246_106# a_381_n377# 0.60fF
C405 s0 a_290_29# 0.60fF
C406 w_738_n73# comp_b2 0.19fF
C407 w_518_405# a_476_404# 2.17fF
C408 a_246_106# a_386_n125# 0.60fF
C409 w_686_n182# D2 0.93fF
C410 w_466_346# a_476_349# 0.42fF
C411 w_738_n18# a_246_106# 1.86fF
C412 a3 a_565_177# 0.87fF
C413 w_561_n319# and_a2 2.64fF
C414 w_613_n411# and_oper_out0 0.19fF
C415 a2 a_565_122# 1.06fF
C416 a_246_106# a_386_n79# 0.60fF
C417 a3 a2 0.41fF
C418 w_332_30# a_246_106# 1.86fF
C419 w_332_30# a_290_29# 2.17fF
C420 a_437_308# b2 0.07fF
C421 a_246_106# a_571_n316# 0.41fF
C422 D1 a_491_234# 0.07fF
C423 a2 D2 0.16fF
C424 a_381_n436# Gnd 6.54fF
C425 and_oper_out0 Gnd 0.88fF
C426 and_b0 Gnd 14.47fF
C427 a_571_n412# Gnd 6.54fF
C428 and_oper_out1 Gnd 0.88fF
C429 a_381_n377# Gnd 6.54fF
C430 and_b1 Gnd 29.42fF
C431 a_571_n360# Gnd 6.54fF
C432 and_oper_out2 Gnd 0.88fF
C433 a_571_n316# Gnd 6.40fF
C434 and_b2 Gnd 28.68fF
C435 a_381_n331# Gnd 6.54fF
C436 and_oper_out3 Gnd 0.88fF
C437 comp_b0 Gnd 0.88fF
C438 a_696_n179# Gnd 6.54fF
C439 a_571_n263# Gnd 6.40fF
C440 comp_b1 Gnd 0.88fF
C441 a_696_n120# Gnd 6.54fF
C442 comp_b2 Gnd 0.88fF
C443 a_696_n74# Gnd 6.54fF
C444 comp_b3 Gnd 0.88fF
C445 a_696_n19# Gnd 6.54fF
C446 comp_a0 Gnd 0.88fF
C447 a_565_17# Gnd 6.54fF
C448 and_b3 Gnd 20.94fF
C449 a_381_n276# Gnd 6.54fF
C450 and_a0 Gnd 43.83fF
C451 a0 Gnd 172.78fF
C452 a_386_n184# Gnd 6.54fF
C453 and_a1 Gnd 12.30fF
C454 a_386_n125# Gnd 6.54fF
C455 and_a2 Gnd 55.92fF
C456 a_386_n79# Gnd 6.54fF
C457 and_a3 Gnd 72.45fF
C458 a_386_n24# Gnd 6.54fF
C459 D3 Gnd 125.71fF
C460 a_290_29# Gnd 6.54fF
C461 comp_a1 Gnd 0.88fF
C462 a_565_76# Gnd 6.54fF
C463 s1 Gnd 35.20fF
C464 a_290_75# Gnd 6.54fF
C465 comp_a2 Gnd 0.88fF
C466 a_565_122# Gnd 6.54fF
C467 comp_a3 Gnd 0.88fF
C468 D2 Gnd 191.11fF
C469 a_565_177# Gnd 6.54fF
C470 adsub_a0 Gnd 0.88fF
C471 a_491_234# Gnd 14.43fF
C472 a_476_244# Gnd 6.54fF
C473 adsub_a1 Gnd 0.88fF
C474 a1 Gnd 38.83fF
C475 a_476_303# Gnd 6.54fF
C476 a_290_124# Gnd 6.54fF
C477 s0 Gnd 61.18fF
C478 s1_not Gnd 11.67fF
C479 s0_not Gnd 21.80fF
C480 a_290_176# Gnd 6.54fF
C481 a_413_308# Gnd 3.59fF
C482 D1 Gnd 51.82fF
C483 D0 Gnd 51.08fF
C484 adsub_a2 Gnd 0.88fF
C485 a2 Gnd 95.62fF
C486 a_476_349# Gnd 6.54fF
C487 adsub_a3 Gnd 0.88fF
C488 a3 Gnd 24.20fF
C489 a_476_404# Gnd 6.54fF
C490 adsub_b0 Gnd 0.88fF
C491 b0 Gnd 320.40fF
C492 a_476_515# Gnd 6.54fF
C493 adsub_b1 Gnd 0.88fF
C494 b1 Gnd 72.08fF
C495 a_476_574# Gnd 6.54fF
C496 adsub_b2 Gnd 0.88fF
C497 b2 Gnd 322.86fF
C498 a_476_620# Gnd 6.54fF
C499 a_246_95# Gnd 370.58fF
C500 adsub_b3 Gnd 0.88fF
C501 a_246_106# Gnd 336.63fF
C502 b3 Gnd 130.59fF
C503 a_437_308# Gnd 115.42fF
C504 a_476_675# Gnd 6.54fF
C505 w_371_n439# Gnd 29.29fF
C506 w_423_n435# Gnd 28.07fF
C507 w_561_n415# Gnd 29.29fF
C508 w_613_n411# Gnd 28.07fF
C509 w_371_n380# Gnd 29.29fF
C510 w_561_n363# Gnd 29.29fF
C511 w_423_n376# Gnd 28.07fF
C512 w_613_n359# Gnd 28.07fF
C513 w_561_n319# Gnd 29.29fF
C514 w_371_n334# Gnd 29.29fF
C515 w_423_n330# Gnd 28.07fF
C516 w_613_n315# Gnd 28.07fF
C517 w_561_n266# Gnd 29.29fF
C518 w_371_n279# Gnd 29.29fF
C519 w_423_n275# Gnd 28.07fF
C520 w_613_n262# Gnd 28.07fF
C521 w_686_n182# Gnd 29.29fF
C522 w_376_n187# Gnd 29.29fF
C523 w_738_n178# Gnd 28.07fF
C524 w_428_n183# Gnd 28.07fF
C525 w_686_n123# Gnd 29.29fF
C526 w_376_n128# Gnd 29.29fF
C527 w_738_n119# Gnd 28.07fF
C528 w_428_n124# Gnd 28.07fF
C529 w_686_n77# Gnd 29.29fF
C530 w_376_n82# Gnd 29.29fF
C531 w_738_n73# Gnd 28.07fF
C532 w_428_n78# Gnd 28.07fF
C533 w_686_n22# Gnd 29.29fF
C534 w_376_n27# Gnd 29.29fF
C535 w_738_n18# Gnd 28.07fF
C536 w_428_n23# Gnd 28.07fF
C537 w_555_14# Gnd 29.29fF
C538 w_607_18# Gnd 28.07fF
C539 w_280_26# Gnd 29.29fF
C540 w_332_30# Gnd 28.07fF
C541 w_555_73# Gnd 29.29fF
C542 w_280_72# Gnd 29.29fF
C543 w_244_81# Gnd 26.36fF
C544 w_607_77# Gnd 28.07fF
C545 w_332_76# Gnd 27.58fF
C546 w_555_119# Gnd 29.29fF
C547 w_607_123# Gnd 28.07fF
C548 w_280_121# Gnd 29.29fF
C549 w_243_117# Gnd 24.41fF
C550 w_332_125# Gnd 27.58fF
C551 w_555_174# Gnd 29.29fF
C552 w_280_173# Gnd 29.29fF
C553 w_607_178# Gnd 28.07fF
C554 w_332_177# Gnd 27.58fF
C555 w_466_241# Gnd 29.29fF
C556 w_518_245# Gnd 28.07fF
C557 w_466_300# Gnd 29.29fF
C558 w_518_304# Gnd 28.07fF
C559 w_404_319# Gnd 41.25fF
C560 w_466_346# Gnd 29.29fF
C561 w_518_350# Gnd 28.07fF
C562 w_466_401# Gnd 29.29fF
C563 w_518_405# Gnd 28.07fF
C564 w_466_512# Gnd 29.29fF
C565 w_518_516# Gnd 28.07fF
C566 w_466_571# Gnd 29.29fF
C567 w_518_575# Gnd 28.07fF
C568 w_466_617# Gnd 29.29fF
C569 w_518_621# Gnd 28.07fF
C570 w_466_672# Gnd 29.29fF
C571 w_518_676# Gnd 28.07fF


.tran 0.1n 800n

.control
run 
* plot v(s0) v(s1)+2
* plot v(D0) v(D1)+2 v(D2)+4 v(D3)+6
plot v(a0) v(a1)+2 v(a2)+4 v(a3)+6
plot v(b0) v(b1)+2 v(b2)+4 v(b3)+6

plot v(and_a0) v(and_a1)+2 v(and_a2)+4 v(and_a3)+6
plot v(and_b0) v(and_b1)+2 v(and_b2)+4 v(and_b3)+6

* plot v(comp_a0) v(comp_a1)+2 v(comp_a2)+4 v(comp_a3)+6
* plot v(comp_b0) v(comp_b1)+2 v(comp_b2)+4 v(comp_b3)+6

* plot v(adsub_a0) v(adsub_a1)+2 v(adsub_a2)+4 v(adsub_a3)+6
* plot v(adsub_b0) v(adsub_b1)+2 v(adsub_b2)+4 v(adsub_b3)+6

* plot v(and_oper_out0) v(and_oper_out1)+2 v(and_oper_out2)+4 v(and_oper_out3)+6
.endc
.endc