magic
tech scmos
timestamp 1700468877
<< nwell >>
rect 477 576 666 630
rect 9 423 333 513
rect 477 468 630 576
rect 477 459 540 468
rect 558 459 630 468
rect 477 99 666 153
rect 9 -54 333 36
rect 477 -9 630 99
rect 477 -18 540 -9
rect 558 -18 630 -9
rect 477 -297 666 -243
rect 9 -450 333 -360
rect 477 -405 630 -297
rect 477 -414 540 -405
rect 558 -414 630 -405
rect 477 -765 666 -711
rect 9 -918 333 -828
rect 477 -873 630 -765
rect 477 -882 540 -873
rect 558 -882 630 -873
<< ntransistor >>
rect 540 378 558 405
rect 81 324 99 351
rect 243 324 261 351
rect 540 -99 558 -72
rect 81 -153 99 -126
rect 243 -153 261 -126
rect 540 -495 558 -468
rect 81 -549 99 -522
rect 243 -549 261 -522
rect 540 -963 558 -936
rect 81 -1017 99 -990
rect 243 -1017 261 -990
<< ptransistor >>
rect 81 450 99 495
rect 243 450 261 495
rect 540 477 558 531
rect 81 -27 99 18
rect 243 -27 261 18
rect 540 0 558 54
rect 81 -423 99 -378
rect 243 -423 261 -378
rect 540 -396 558 -342
rect 81 -891 99 -846
rect 243 -891 261 -846
rect 540 -864 558 -810
<< ndiffusion >>
rect 495 396 540 405
rect 495 378 504 396
rect 531 378 540 396
rect 558 378 576 405
rect 603 378 612 405
rect 45 342 81 351
rect 45 324 54 342
rect 72 324 81 342
rect 99 324 243 351
rect 261 333 270 351
rect 288 333 297 351
rect 261 324 297 333
rect 495 -81 540 -72
rect 495 -99 504 -81
rect 531 -99 540 -81
rect 558 -99 576 -72
rect 603 -99 612 -72
rect 45 -135 81 -126
rect 45 -153 54 -135
rect 72 -153 81 -135
rect 99 -153 243 -126
rect 261 -144 270 -126
rect 288 -144 297 -126
rect 261 -153 297 -144
rect 495 -477 540 -468
rect 495 -495 504 -477
rect 531 -495 540 -477
rect 558 -495 576 -468
rect 603 -495 612 -468
rect 45 -531 81 -522
rect 45 -549 54 -531
rect 72 -549 81 -531
rect 99 -549 243 -522
rect 261 -540 270 -522
rect 288 -540 297 -522
rect 261 -549 297 -540
rect 495 -945 540 -936
rect 495 -963 504 -945
rect 531 -963 540 -945
rect 558 -963 576 -936
rect 603 -963 612 -936
rect 45 -999 81 -990
rect 45 -1017 54 -999
rect 72 -1017 81 -999
rect 99 -1017 243 -990
rect 261 -1008 270 -990
rect 288 -1008 297 -990
rect 261 -1017 297 -1008
<< pdiffusion >>
rect 495 504 504 531
rect 531 504 540 531
rect 45 486 81 495
rect 45 468 54 486
rect 72 468 81 486
rect 45 450 81 468
rect 99 477 162 495
rect 99 459 108 477
rect 126 459 162 477
rect 99 450 162 459
rect 198 486 243 495
rect 198 468 207 486
rect 225 468 243 486
rect 198 450 243 468
rect 261 486 297 495
rect 261 468 270 486
rect 288 468 297 486
rect 495 477 540 504
rect 558 522 612 531
rect 558 495 576 522
rect 603 495 612 522
rect 558 477 612 495
rect 261 450 297 468
rect 495 27 504 54
rect 531 27 540 54
rect 45 9 81 18
rect 45 -9 54 9
rect 72 -9 81 9
rect 45 -27 81 -9
rect 99 0 162 18
rect 99 -18 108 0
rect 126 -18 162 0
rect 99 -27 162 -18
rect 198 9 243 18
rect 198 -9 207 9
rect 225 -9 243 9
rect 198 -27 243 -9
rect 261 9 297 18
rect 261 -9 270 9
rect 288 -9 297 9
rect 495 0 540 27
rect 558 45 612 54
rect 558 18 576 45
rect 603 18 612 45
rect 558 0 612 18
rect 261 -27 297 -9
rect 495 -369 504 -342
rect 531 -369 540 -342
rect 45 -387 81 -378
rect 45 -405 54 -387
rect 72 -405 81 -387
rect 45 -423 81 -405
rect 99 -396 162 -378
rect 99 -414 108 -396
rect 126 -414 162 -396
rect 99 -423 162 -414
rect 198 -387 243 -378
rect 198 -405 207 -387
rect 225 -405 243 -387
rect 198 -423 243 -405
rect 261 -387 297 -378
rect 261 -405 270 -387
rect 288 -405 297 -387
rect 495 -396 540 -369
rect 558 -351 612 -342
rect 558 -378 576 -351
rect 603 -378 612 -351
rect 558 -396 612 -378
rect 261 -423 297 -405
rect 495 -837 504 -810
rect 531 -837 540 -810
rect 45 -855 81 -846
rect 45 -873 54 -855
rect 72 -873 81 -855
rect 45 -891 81 -873
rect 99 -864 162 -846
rect 99 -882 108 -864
rect 126 -882 162 -864
rect 99 -891 162 -882
rect 198 -855 243 -846
rect 198 -873 207 -855
rect 225 -873 243 -855
rect 198 -891 243 -873
rect 261 -855 297 -846
rect 261 -873 270 -855
rect 288 -873 297 -855
rect 495 -864 540 -837
rect 558 -819 612 -810
rect 558 -846 576 -819
rect 603 -846 612 -819
rect 558 -864 612 -846
rect 261 -891 297 -873
<< ndcontact >>
rect 504 369 531 396
rect 576 378 603 405
rect 54 324 72 342
rect 270 333 288 351
rect 504 -108 531 -81
rect 576 -99 603 -72
rect 54 -153 72 -135
rect 270 -144 288 -126
rect 504 -504 531 -477
rect 576 -495 603 -468
rect 54 -549 72 -531
rect 270 -540 288 -522
rect 504 -972 531 -945
rect 576 -963 603 -936
rect 54 -1017 72 -999
rect 270 -1008 288 -990
<< pdcontact >>
rect 504 504 531 531
rect 54 468 72 486
rect 108 459 126 477
rect 207 468 225 486
rect 270 468 288 486
rect 576 495 603 522
rect 504 27 531 54
rect 54 -9 72 9
rect 108 -18 126 0
rect 207 -9 225 9
rect 270 -9 288 9
rect 576 18 603 45
rect 504 -369 531 -342
rect 54 -405 72 -387
rect 108 -414 126 -396
rect 207 -405 225 -387
rect 270 -405 288 -387
rect 576 -378 603 -351
rect 504 -837 531 -810
rect 54 -873 72 -855
rect 108 -882 126 -864
rect 207 -873 225 -855
rect 270 -873 288 -855
rect 576 -846 603 -819
<< polysilicon >>
rect 540 531 558 648
rect 81 495 99 522
rect 243 495 261 522
rect 81 351 99 450
rect 243 351 261 450
rect 540 441 558 477
rect 549 414 558 441
rect 540 405 558 414
rect 540 360 558 378
rect 81 315 99 324
rect 243 315 261 324
rect 540 54 558 171
rect 81 18 99 45
rect 243 18 261 45
rect 81 -126 99 -27
rect 243 -126 261 -27
rect 540 -36 558 0
rect 549 -63 558 -36
rect 540 -72 558 -63
rect 540 -117 558 -99
rect 81 -162 99 -153
rect 243 -162 261 -153
rect 540 -342 558 -225
rect 81 -378 99 -351
rect 243 -378 261 -351
rect 81 -522 99 -423
rect 243 -522 261 -423
rect 540 -432 558 -396
rect 549 -459 558 -432
rect 540 -468 558 -459
rect 540 -513 558 -495
rect 81 -558 99 -549
rect 243 -558 261 -549
rect 540 -810 558 -693
rect 81 -846 99 -819
rect 243 -846 261 -819
rect 81 -990 99 -891
rect 243 -990 261 -891
rect 540 -900 558 -864
rect 549 -927 558 -900
rect 540 -936 558 -927
rect 540 -981 558 -963
rect 81 -1026 99 -1017
rect 243 -1026 261 -1017
<< polycontact >>
rect 522 414 549 441
rect 522 -63 549 -36
rect 522 -459 549 -432
rect 522 -927 549 -900
<< metal1 >>
rect 504 585 603 594
rect 504 558 531 585
rect -108 540 531 558
rect -108 81 -90 540
rect 54 486 72 540
rect 207 486 225 540
rect 504 531 531 540
rect 108 405 126 459
rect 270 405 288 468
rect 576 450 603 495
rect 432 414 522 441
rect 576 423 630 450
rect 432 405 450 414
rect 108 387 450 405
rect 576 405 603 423
rect 270 351 288 387
rect 504 342 531 369
rect 54 306 72 324
rect 504 324 720 342
rect 504 306 540 324
rect 54 288 540 306
rect 504 108 603 117
rect 504 81 531 108
rect -108 63 531 81
rect -108 -315 -90 63
rect 54 9 72 63
rect 207 9 225 63
rect 504 54 531 63
rect 108 -72 126 -18
rect 270 -72 288 -9
rect 576 -27 603 18
rect 432 -63 522 -36
rect 576 -54 630 -27
rect 432 -72 450 -63
rect 108 -90 450 -72
rect 576 -72 603 -54
rect 270 -126 288 -90
rect 504 -135 531 -108
rect 702 -135 720 324
rect 54 -171 72 -153
rect 504 -153 720 -135
rect 504 -171 540 -153
rect 54 -189 540 -171
rect 504 -288 603 -279
rect 504 -315 531 -288
rect -108 -333 531 -315
rect -108 -783 -90 -333
rect 54 -387 72 -333
rect 207 -387 225 -333
rect 504 -342 531 -333
rect 108 -468 126 -414
rect 270 -468 288 -405
rect 576 -423 603 -378
rect 432 -459 522 -432
rect 576 -450 630 -423
rect 432 -468 450 -459
rect 108 -486 450 -468
rect 576 -468 603 -450
rect 270 -522 288 -486
rect 504 -531 531 -504
rect 702 -531 720 -153
rect 54 -567 72 -549
rect 504 -549 720 -531
rect 504 -567 540 -549
rect 54 -585 540 -567
rect 504 -756 603 -747
rect 504 -783 531 -756
rect -108 -801 531 -783
rect 54 -855 72 -801
rect 207 -855 225 -801
rect 504 -810 531 -801
rect 108 -936 126 -882
rect 270 -936 288 -873
rect 576 -891 603 -846
rect 432 -927 522 -900
rect 576 -918 630 -891
rect 432 -936 450 -927
rect 108 -954 450 -936
rect 576 -936 603 -918
rect 270 -990 288 -954
rect 504 -999 531 -972
rect 702 -999 720 -549
rect 54 -1035 72 -1017
rect 504 -1017 720 -999
rect 504 -1035 540 -1017
rect 54 -1053 540 -1035
<< labels >>
rlabel polysilicon 90 -945 90 -945 1 a0
rlabel polysilicon 252 -963 252 -963 1 b0
rlabel metal1 603 -900 603 -900 1 and_oper_out0
rlabel polysilicon 90 -477 90 -477 1 a1
rlabel polysilicon 252 -504 252 -504 1 b1
rlabel metal1 603 -432 603 -432 1 and_oper_out1
rlabel polysilicon 90 -108 90 -108 1 a2
rlabel polysilicon 252 -108 252 -108 1 b2
rlabel metal1 612 -45 612 -45 1 and_oper_out2
rlabel polysilicon 90 378 90 378 1 a3
rlabel polysilicon 252 369 252 369 1 b3
rlabel metal1 612 432 612 432 1 and_oper_out3
rlabel metal1 288 -576 288 -576 1 gnd
rlabel metal1 -81 -324 -81 -324 3 vdd
<< end >>
