magic
tech scmos
magscale 9 1
timestamp 1700391575
<< nwell >>
rect -10 10 11 15
rect -9 -2 8 10
rect -9 -3 -2 -2
rect 0 -3 8 -2
<< ntransistor >>
rect -2 -12 0 -9
<< ptransistor >>
rect -2 -1 0 5
<< ndiffusion >>
rect -7 -10 -2 -9
rect -7 -12 -6 -10
rect -3 -12 -2 -10
rect 0 -12 2 -9
rect 5 -12 6 -9
<< pdiffusion >>
rect -7 2 -6 5
rect -3 2 -2 5
rect -7 -1 -2 2
rect 0 4 6 5
rect 0 1 2 4
rect 5 1 6 4
rect 0 -1 6 1
<< ndcontact >>
rect -6 -13 -3 -10
rect 2 -12 5 -9
<< pdcontact >>
rect -6 2 -3 5
rect 2 1 5 4
<< polysilicon >>
rect -2 5 0 7
rect -2 -5 0 -1
rect -1 -8 0 -5
rect -2 -9 0 -8
rect -2 -14 0 -12
<< polycontact >>
rect -4 -8 -1 -5
<< metal1 >>
rect -7 11 5 12
rect -7 10 -3 11
rect -6 5 -3 10
rect 2 -4 5 1
rect -6 -8 -4 -5
rect 2 -7 8 -4
rect 2 -9 5 -7
rect -6 -16 -3 -13
rect -7 -18 4 -16
<< labels >>
rlabel metal1 -6 -7 -6 -7 1 A
rlabel metal1 4 -7 4 -7 1 out
rlabel metal1 -6 11 -6 11 1 vdd
rlabel metal1 -1 -18 -1 -18 1 gnd
<< end >>
