magic
tech scmos
timestamp 1701034540
<< nwell >>
rect 4554 4797 4743 4851
rect 4086 4644 4410 4734
rect 4554 4689 4707 4797
rect 4554 4680 4617 4689
rect 4635 4680 4707 4689
rect 4554 4302 4743 4356
rect 4086 4149 4410 4239
rect 4554 4194 4707 4302
rect 4554 4185 4617 4194
rect 4635 4185 4707 4194
rect 3528 3906 3879 4023
rect 4554 3888 4743 3942
rect 4086 3735 4410 3825
rect 4554 3780 4707 3888
rect 4554 3771 4617 3780
rect 4635 3771 4707 3780
rect 4554 3357 4743 3411
rect 4086 3204 4410 3294
rect 4554 3249 4707 3357
rect 4554 3240 4617 3249
rect 4635 3240 4707 3249
rect 4554 2790 4743 2844
rect 4086 2637 4410 2727
rect 4554 2682 4707 2790
rect 4554 2673 4617 2682
rect 4635 2673 4707 2682
rect 4554 2295 4743 2349
rect 4086 2142 4410 2232
rect 4554 2187 4707 2295
rect 4554 2178 4617 2187
rect 4635 2178 4707 2187
rect 4554 1881 4743 1935
rect 4086 1728 4410 1818
rect 4554 1773 4707 1881
rect 4554 1764 4617 1773
rect 4635 1764 4707 1773
rect 2601 1674 2790 1728
rect 2133 1521 2457 1611
rect 2601 1566 2754 1674
rect 2601 1557 2664 1566
rect 2682 1557 2754 1566
rect 4554 1350 4743 1404
rect 2601 1206 2790 1260
rect 1800 1035 1989 1062
rect 2133 1053 2457 1143
rect 2601 1098 2754 1206
rect 4086 1197 4410 1287
rect 4554 1242 4707 1350
rect 4554 1233 4617 1242
rect 4635 1233 4707 1242
rect 2601 1089 2664 1098
rect 2682 1089 2754 1098
rect 1800 1017 1827 1035
rect 1935 1017 1989 1035
rect 1809 909 1962 1017
rect 1809 900 1872 909
rect 1890 900 1962 909
rect 2601 765 2790 819
rect 4545 801 4734 855
rect 1809 720 1998 738
rect 2070 720 2088 747
rect 1809 702 2088 720
rect 1809 693 1998 702
rect 1818 585 1971 693
rect 2133 612 2457 702
rect 2601 657 2754 765
rect 2601 648 2664 657
rect 2682 648 2754 657
rect 4077 648 4401 738
rect 4545 693 4698 801
rect 4545 684 4608 693
rect 4626 684 4698 693
rect 1818 576 1881 585
rect 1899 576 1971 585
rect 2601 351 2790 405
rect 2133 198 2457 288
rect 2601 243 2754 351
rect 4545 306 4734 360
rect 2601 234 2664 243
rect 2682 234 2754 243
rect 4077 153 4401 243
rect 4545 198 4698 306
rect 4545 189 4608 198
rect 4626 189 4698 198
rect 4545 -108 4734 -54
rect 4077 -261 4401 -171
rect 4545 -216 4698 -108
rect 4545 -225 4608 -216
rect 4626 -225 4698 -216
rect 4545 -639 4734 -585
rect 4077 -792 4401 -702
rect 4545 -747 4698 -639
rect 4545 -756 4608 -747
rect 4626 -756 4698 -747
rect 4545 -1116 4734 -1062
rect 4077 -1269 4401 -1179
rect 4545 -1224 4698 -1116
rect 4545 -1233 4608 -1224
rect 4626 -1233 4698 -1224
rect 4545 -1611 4734 -1557
rect 4077 -1764 4401 -1674
rect 4545 -1719 4698 -1611
rect 4545 -1728 4608 -1719
rect 4626 -1728 4698 -1719
rect 4545 -2025 4734 -1971
rect 4077 -2178 4401 -2088
rect 4545 -2133 4698 -2025
rect 4545 -2142 4608 -2133
rect 4626 -2142 4698 -2133
rect 4545 -2556 4734 -2502
rect 4077 -2709 4401 -2619
rect 4545 -2664 4698 -2556
rect 4545 -2673 4608 -2664
rect 4626 -2673 4698 -2664
rect 4545 -3123 4734 -3069
rect 4077 -3276 4401 -3186
rect 4545 -3231 4698 -3123
rect 4545 -3240 4608 -3231
rect 4626 -3240 4698 -3231
rect 4545 -3618 4734 -3564
rect 4077 -3771 4401 -3681
rect 4545 -3726 4698 -3618
rect 4545 -3735 4608 -3726
rect 4626 -3735 4698 -3726
rect 4545 -4032 4734 -3978
rect 4077 -4185 4401 -4095
rect 4545 -4140 4698 -4032
rect 4545 -4149 4608 -4140
rect 4626 -4149 4698 -4140
rect 4545 -4563 4734 -4509
rect 4077 -4716 4401 -4626
rect 4545 -4671 4698 -4563
rect 4545 -4680 4608 -4671
rect 4626 -4680 4698 -4671
rect 4545 -5058 4734 -5004
rect 4077 -5211 4401 -5121
rect 4545 -5166 4698 -5058
rect 4545 -5175 4608 -5166
rect 4626 -5175 4698 -5166
rect 4545 -5553 4734 -5499
rect 4077 -5706 4401 -5616
rect 4545 -5661 4698 -5553
rect 4545 -5670 4608 -5661
rect 4626 -5670 4698 -5661
rect 4545 -5967 4734 -5913
rect 4077 -6120 4401 -6030
rect 4545 -6075 4698 -5967
rect 4545 -6084 4608 -6075
rect 4626 -6084 4698 -6075
rect 4545 -6498 4734 -6444
rect 4077 -6651 4401 -6561
rect 4545 -6606 4698 -6498
rect 4545 -6615 4608 -6606
rect 4626 -6615 4698 -6606
<< ntransistor >>
rect 4617 4599 4635 4626
rect 4158 4545 4176 4572
rect 4320 4545 4338 4572
rect 4617 4104 4635 4131
rect 4158 4050 4176 4077
rect 4320 4050 4338 4077
rect 3591 3807 3609 3834
rect 3681 3807 3699 3834
rect 3807 3807 3825 3834
rect 2664 1476 2682 1503
rect 2205 1422 2223 1449
rect 2367 1422 2385 1449
rect 4617 3690 4635 3717
rect 4158 3636 4176 3663
rect 4320 3636 4338 3663
rect 4617 3159 4635 3186
rect 4158 3105 4176 3132
rect 4320 3105 4338 3132
rect 4617 2592 4635 2619
rect 4158 2538 4176 2565
rect 4320 2538 4338 2565
rect 4617 2097 4635 2124
rect 4158 2043 4176 2070
rect 4320 2043 4338 2070
rect 4617 1683 4635 1710
rect 4158 1629 4176 1656
rect 4320 1629 4338 1656
rect 4617 1152 4635 1179
rect 4158 1098 4176 1125
rect 4320 1098 4338 1125
rect 2664 1008 2682 1035
rect 2205 954 2223 981
rect 2367 954 2385 981
rect 1872 819 1890 846
rect 2664 567 2682 594
rect 1881 495 1899 522
rect 2205 513 2223 540
rect 2340 513 2358 540
rect 2367 513 2385 540
rect 2664 153 2682 180
rect 2205 99 2223 126
rect 2322 99 2340 126
rect 2367 99 2385 126
rect 4608 603 4626 630
rect 4149 549 4167 576
rect 4311 549 4329 576
rect 4608 108 4626 135
rect 4149 54 4167 81
rect 4311 54 4329 81
rect 4608 -306 4626 -279
rect 4149 -360 4167 -333
rect 4311 -360 4329 -333
rect 4608 -837 4626 -810
rect 4149 -891 4167 -864
rect 4311 -891 4329 -864
rect 4608 -1314 4626 -1287
rect 4149 -1368 4167 -1341
rect 4311 -1368 4329 -1341
rect 4608 -1809 4626 -1782
rect 4149 -1863 4167 -1836
rect 4311 -1863 4329 -1836
rect 4608 -2223 4626 -2196
rect 4149 -2277 4167 -2250
rect 4311 -2277 4329 -2250
rect 4608 -2754 4626 -2727
rect 4149 -2808 4167 -2781
rect 4311 -2808 4329 -2781
rect 4608 -3321 4626 -3294
rect 4149 -3375 4167 -3348
rect 4311 -3375 4329 -3348
rect 4608 -3816 4626 -3789
rect 4149 -3870 4167 -3843
rect 4311 -3870 4329 -3843
rect 4608 -4230 4626 -4203
rect 4149 -4284 4167 -4257
rect 4311 -4284 4329 -4257
rect 4608 -4761 4626 -4734
rect 4149 -4815 4167 -4788
rect 4311 -4815 4329 -4788
rect 4608 -5256 4626 -5229
rect 4149 -5310 4167 -5283
rect 4311 -5310 4329 -5283
rect 4608 -5751 4626 -5724
rect 4149 -5805 4167 -5778
rect 4311 -5805 4329 -5778
rect 4608 -6165 4626 -6138
rect 4149 -6219 4167 -6192
rect 4311 -6219 4329 -6192
rect 4608 -6696 4626 -6669
rect 4149 -6750 4167 -6723
rect 4311 -6750 4329 -6723
<< ptransistor >>
rect 4158 4671 4176 4716
rect 4320 4671 4338 4716
rect 4617 4698 4635 4752
rect 4158 4176 4176 4221
rect 4320 4176 4338 4221
rect 4617 4203 4635 4257
rect 3591 3924 3609 3969
rect 3681 3924 3699 3969
rect 3807 3924 3825 3969
rect 2205 1548 2223 1593
rect 2367 1548 2385 1593
rect 2664 1575 2682 1629
rect 4158 3762 4176 3807
rect 4320 3762 4338 3807
rect 4617 3789 4635 3843
rect 2205 1080 2223 1125
rect 2367 1080 2385 1125
rect 2664 1107 2682 1161
rect 4158 3231 4176 3276
rect 4320 3231 4338 3276
rect 4617 3258 4635 3312
rect 4158 2664 4176 2709
rect 4320 2664 4338 2709
rect 4617 2691 4635 2745
rect 4158 2169 4176 2214
rect 4320 2169 4338 2214
rect 4617 2196 4635 2250
rect 4158 1755 4176 1800
rect 4320 1755 4338 1800
rect 4617 1782 4635 1836
rect 4158 1224 4176 1269
rect 4320 1224 4338 1269
rect 4617 1251 4635 1305
rect 1872 918 1890 972
rect 1881 594 1899 648
rect 2205 639 2223 684
rect 2367 639 2385 684
rect 2664 666 2682 720
rect 4149 675 4167 720
rect 4311 675 4329 720
rect 4608 702 4626 756
rect 2205 225 2223 270
rect 2367 225 2385 270
rect 2664 252 2682 306
rect 4149 180 4167 225
rect 4311 180 4329 225
rect 4608 207 4626 261
rect 4149 -234 4167 -189
rect 4311 -234 4329 -189
rect 4608 -207 4626 -153
rect 4149 -765 4167 -720
rect 4311 -765 4329 -720
rect 4608 -738 4626 -684
rect 4149 -1242 4167 -1197
rect 4311 -1242 4329 -1197
rect 4608 -1215 4626 -1161
rect 4149 -1737 4167 -1692
rect 4311 -1737 4329 -1692
rect 4608 -1710 4626 -1656
rect 4149 -2151 4167 -2106
rect 4311 -2151 4329 -2106
rect 4608 -2124 4626 -2070
rect 4149 -2682 4167 -2637
rect 4311 -2682 4329 -2637
rect 4608 -2655 4626 -2601
rect 4149 -3249 4167 -3204
rect 4311 -3249 4329 -3204
rect 4608 -3222 4626 -3168
rect 4149 -3744 4167 -3699
rect 4311 -3744 4329 -3699
rect 4608 -3717 4626 -3663
rect 4149 -4158 4167 -4113
rect 4311 -4158 4329 -4113
rect 4608 -4131 4626 -4077
rect 4149 -4689 4167 -4644
rect 4311 -4689 4329 -4644
rect 4608 -4662 4626 -4608
rect 4149 -5184 4167 -5139
rect 4311 -5184 4329 -5139
rect 4608 -5157 4626 -5103
rect 4149 -5679 4167 -5634
rect 4311 -5679 4329 -5634
rect 4608 -5652 4626 -5598
rect 4149 -6093 4167 -6048
rect 4311 -6093 4329 -6048
rect 4608 -6066 4626 -6012
rect 4149 -6624 4167 -6579
rect 4311 -6624 4329 -6579
rect 4608 -6597 4626 -6543
<< ndiffusion >>
rect 4572 4617 4617 4626
rect 4572 4599 4581 4617
rect 4608 4599 4617 4617
rect 4635 4599 4653 4626
rect 4680 4599 4689 4626
rect 4122 4563 4158 4572
rect 4122 4545 4131 4563
rect 4149 4545 4158 4563
rect 4176 4545 4320 4572
rect 4338 4554 4347 4572
rect 4365 4554 4374 4572
rect 4338 4545 4374 4554
rect 4572 4122 4617 4131
rect 4572 4104 4581 4122
rect 4608 4104 4617 4122
rect 4635 4104 4653 4131
rect 4680 4104 4689 4131
rect 4122 4068 4158 4077
rect 4122 4050 4131 4068
rect 4149 4050 4158 4068
rect 4176 4050 4320 4077
rect 4338 4059 4347 4077
rect 4365 4059 4374 4077
rect 4338 4050 4374 4059
rect 3555 3816 3564 3834
rect 3582 3816 3591 3834
rect 3555 3807 3591 3816
rect 3609 3816 3618 3834
rect 3609 3807 3636 3816
rect 3645 3816 3654 3834
rect 3672 3816 3681 3834
rect 3645 3807 3681 3816
rect 3699 3816 3708 3834
rect 3699 3807 3726 3816
rect 3771 3816 3780 3834
rect 3798 3816 3807 3834
rect 3771 3807 3807 3816
rect 3825 3816 3834 3834
rect 3852 3816 3861 3834
rect 3825 3807 3861 3816
rect 2619 1494 2664 1503
rect 2619 1476 2628 1494
rect 2655 1476 2664 1494
rect 2682 1476 2700 1503
rect 2727 1476 2736 1503
rect 2169 1440 2205 1449
rect 2169 1422 2178 1440
rect 2196 1422 2205 1440
rect 2223 1422 2367 1449
rect 2385 1431 2394 1449
rect 2412 1431 2421 1449
rect 2385 1422 2421 1431
rect 4572 3708 4617 3717
rect 4572 3690 4581 3708
rect 4608 3690 4617 3708
rect 4635 3690 4653 3717
rect 4680 3690 4689 3717
rect 4122 3654 4158 3663
rect 4122 3636 4131 3654
rect 4149 3636 4158 3654
rect 4176 3636 4320 3663
rect 4338 3645 4347 3663
rect 4365 3645 4374 3663
rect 4338 3636 4374 3645
rect 4572 3177 4617 3186
rect 4572 3159 4581 3177
rect 4608 3159 4617 3177
rect 4635 3159 4653 3186
rect 4680 3159 4689 3186
rect 4122 3123 4158 3132
rect 4122 3105 4131 3123
rect 4149 3105 4158 3123
rect 4176 3105 4320 3132
rect 4338 3114 4347 3132
rect 4365 3114 4374 3132
rect 4338 3105 4374 3114
rect 4572 2610 4617 2619
rect 4572 2592 4581 2610
rect 4608 2592 4617 2610
rect 4635 2592 4653 2619
rect 4680 2592 4689 2619
rect 4122 2556 4158 2565
rect 4122 2538 4131 2556
rect 4149 2538 4158 2556
rect 4176 2538 4320 2565
rect 4338 2547 4347 2565
rect 4365 2547 4374 2565
rect 4338 2538 4374 2547
rect 4572 2115 4617 2124
rect 4572 2097 4581 2115
rect 4608 2097 4617 2115
rect 4635 2097 4653 2124
rect 4680 2097 4689 2124
rect 4122 2061 4158 2070
rect 4122 2043 4131 2061
rect 4149 2043 4158 2061
rect 4176 2043 4320 2070
rect 4338 2052 4347 2070
rect 4365 2052 4374 2070
rect 4338 2043 4374 2052
rect 4572 1701 4617 1710
rect 4572 1683 4581 1701
rect 4608 1683 4617 1701
rect 4635 1683 4653 1710
rect 4680 1683 4689 1710
rect 4122 1647 4158 1656
rect 4122 1629 4131 1647
rect 4149 1629 4158 1647
rect 4176 1629 4320 1656
rect 4338 1638 4347 1656
rect 4365 1638 4374 1656
rect 4338 1629 4374 1638
rect 4572 1170 4617 1179
rect 4572 1152 4581 1170
rect 4608 1152 4617 1170
rect 4635 1152 4653 1179
rect 4680 1152 4689 1179
rect 4122 1116 4158 1125
rect 4122 1098 4131 1116
rect 4149 1098 4158 1116
rect 4176 1098 4320 1125
rect 4338 1107 4347 1125
rect 4365 1107 4374 1125
rect 4338 1098 4374 1107
rect 2619 1026 2664 1035
rect 2619 1008 2628 1026
rect 2655 1008 2664 1026
rect 2682 1008 2700 1035
rect 2727 1008 2736 1035
rect 2169 972 2205 981
rect 2169 954 2178 972
rect 2196 954 2205 972
rect 2223 954 2367 981
rect 2385 963 2394 981
rect 2412 963 2421 981
rect 2385 954 2421 963
rect 1827 837 1872 846
rect 1827 819 1836 837
rect 1863 819 1872 837
rect 1890 819 1908 846
rect 1935 819 1944 846
rect 2619 585 2664 594
rect 2619 567 2628 585
rect 2655 567 2664 585
rect 2682 567 2700 594
rect 2727 567 2736 594
rect 2169 531 2205 540
rect 1836 513 1881 522
rect 1836 495 1845 513
rect 1872 495 1881 513
rect 1899 495 1917 522
rect 1944 495 1953 522
rect 2169 513 2178 531
rect 2196 513 2205 531
rect 2223 513 2340 540
rect 2358 513 2367 540
rect 2385 522 2394 540
rect 2412 522 2421 540
rect 2385 513 2421 522
rect 2619 171 2664 180
rect 2619 153 2628 171
rect 2655 153 2664 171
rect 2682 153 2700 180
rect 2727 153 2736 180
rect 2169 117 2205 126
rect 2169 99 2178 117
rect 2196 99 2205 117
rect 2223 99 2322 126
rect 2340 99 2367 126
rect 2385 108 2394 126
rect 2412 108 2421 126
rect 2385 99 2421 108
rect 4563 621 4608 630
rect 4563 603 4572 621
rect 4599 603 4608 621
rect 4626 603 4644 630
rect 4671 603 4680 630
rect 4113 567 4149 576
rect 4113 549 4122 567
rect 4140 549 4149 567
rect 4167 549 4311 576
rect 4329 558 4338 576
rect 4356 558 4365 576
rect 4329 549 4365 558
rect 4563 126 4608 135
rect 4563 108 4572 126
rect 4599 108 4608 126
rect 4626 108 4644 135
rect 4671 108 4680 135
rect 4113 72 4149 81
rect 4113 54 4122 72
rect 4140 54 4149 72
rect 4167 54 4311 81
rect 4329 63 4338 81
rect 4356 63 4365 81
rect 4329 54 4365 63
rect 4563 -288 4608 -279
rect 4563 -306 4572 -288
rect 4599 -306 4608 -288
rect 4626 -306 4644 -279
rect 4671 -306 4680 -279
rect 4113 -342 4149 -333
rect 4113 -360 4122 -342
rect 4140 -360 4149 -342
rect 4167 -360 4311 -333
rect 4329 -351 4338 -333
rect 4356 -351 4365 -333
rect 4329 -360 4365 -351
rect 4563 -819 4608 -810
rect 4563 -837 4572 -819
rect 4599 -837 4608 -819
rect 4626 -837 4644 -810
rect 4671 -837 4680 -810
rect 4113 -873 4149 -864
rect 4113 -891 4122 -873
rect 4140 -891 4149 -873
rect 4167 -891 4311 -864
rect 4329 -882 4338 -864
rect 4356 -882 4365 -864
rect 4329 -891 4365 -882
rect 4563 -1296 4608 -1287
rect 4563 -1314 4572 -1296
rect 4599 -1314 4608 -1296
rect 4626 -1314 4644 -1287
rect 4671 -1314 4680 -1287
rect 4113 -1350 4149 -1341
rect 4113 -1368 4122 -1350
rect 4140 -1368 4149 -1350
rect 4167 -1368 4311 -1341
rect 4329 -1359 4338 -1341
rect 4356 -1359 4365 -1341
rect 4329 -1368 4365 -1359
rect 4563 -1791 4608 -1782
rect 4563 -1809 4572 -1791
rect 4599 -1809 4608 -1791
rect 4626 -1809 4644 -1782
rect 4671 -1809 4680 -1782
rect 4113 -1845 4149 -1836
rect 4113 -1863 4122 -1845
rect 4140 -1863 4149 -1845
rect 4167 -1863 4311 -1836
rect 4329 -1854 4338 -1836
rect 4356 -1854 4365 -1836
rect 4329 -1863 4365 -1854
rect 4563 -2205 4608 -2196
rect 4563 -2223 4572 -2205
rect 4599 -2223 4608 -2205
rect 4626 -2223 4644 -2196
rect 4671 -2223 4680 -2196
rect 4113 -2259 4149 -2250
rect 4113 -2277 4122 -2259
rect 4140 -2277 4149 -2259
rect 4167 -2277 4311 -2250
rect 4329 -2268 4338 -2250
rect 4356 -2268 4365 -2250
rect 4329 -2277 4365 -2268
rect 4563 -2736 4608 -2727
rect 4563 -2754 4572 -2736
rect 4599 -2754 4608 -2736
rect 4626 -2754 4644 -2727
rect 4671 -2754 4680 -2727
rect 4113 -2790 4149 -2781
rect 4113 -2808 4122 -2790
rect 4140 -2808 4149 -2790
rect 4167 -2808 4311 -2781
rect 4329 -2799 4338 -2781
rect 4356 -2799 4365 -2781
rect 4329 -2808 4365 -2799
rect 4563 -3303 4608 -3294
rect 4563 -3321 4572 -3303
rect 4599 -3321 4608 -3303
rect 4626 -3321 4644 -3294
rect 4671 -3321 4680 -3294
rect 4113 -3357 4149 -3348
rect 4113 -3375 4122 -3357
rect 4140 -3375 4149 -3357
rect 4167 -3375 4311 -3348
rect 4329 -3366 4338 -3348
rect 4356 -3366 4365 -3348
rect 4329 -3375 4365 -3366
rect 4563 -3798 4608 -3789
rect 4563 -3816 4572 -3798
rect 4599 -3816 4608 -3798
rect 4626 -3816 4644 -3789
rect 4671 -3816 4680 -3789
rect 4113 -3852 4149 -3843
rect 4113 -3870 4122 -3852
rect 4140 -3870 4149 -3852
rect 4167 -3870 4311 -3843
rect 4329 -3861 4338 -3843
rect 4356 -3861 4365 -3843
rect 4329 -3870 4365 -3861
rect 4563 -4212 4608 -4203
rect 4563 -4230 4572 -4212
rect 4599 -4230 4608 -4212
rect 4626 -4230 4644 -4203
rect 4671 -4230 4680 -4203
rect 4113 -4266 4149 -4257
rect 4113 -4284 4122 -4266
rect 4140 -4284 4149 -4266
rect 4167 -4284 4311 -4257
rect 4329 -4275 4338 -4257
rect 4356 -4275 4365 -4257
rect 4329 -4284 4365 -4275
rect 4563 -4743 4608 -4734
rect 4563 -4761 4572 -4743
rect 4599 -4761 4608 -4743
rect 4626 -4761 4644 -4734
rect 4671 -4761 4680 -4734
rect 4113 -4797 4149 -4788
rect 4113 -4815 4122 -4797
rect 4140 -4815 4149 -4797
rect 4167 -4815 4311 -4788
rect 4329 -4806 4338 -4788
rect 4356 -4806 4365 -4788
rect 4329 -4815 4365 -4806
rect 4563 -5238 4608 -5229
rect 4563 -5256 4572 -5238
rect 4599 -5256 4608 -5238
rect 4626 -5256 4644 -5229
rect 4671 -5256 4680 -5229
rect 4113 -5292 4149 -5283
rect 4113 -5310 4122 -5292
rect 4140 -5310 4149 -5292
rect 4167 -5310 4311 -5283
rect 4329 -5301 4338 -5283
rect 4356 -5301 4365 -5283
rect 4329 -5310 4365 -5301
rect 4563 -5733 4608 -5724
rect 4563 -5751 4572 -5733
rect 4599 -5751 4608 -5733
rect 4626 -5751 4644 -5724
rect 4671 -5751 4680 -5724
rect 4113 -5787 4149 -5778
rect 4113 -5805 4122 -5787
rect 4140 -5805 4149 -5787
rect 4167 -5805 4311 -5778
rect 4329 -5796 4338 -5778
rect 4356 -5796 4365 -5778
rect 4329 -5805 4365 -5796
rect 4563 -6147 4608 -6138
rect 4563 -6165 4572 -6147
rect 4599 -6165 4608 -6147
rect 4626 -6165 4644 -6138
rect 4671 -6165 4680 -6138
rect 4113 -6201 4149 -6192
rect 4113 -6219 4122 -6201
rect 4140 -6219 4149 -6201
rect 4167 -6219 4311 -6192
rect 4329 -6210 4338 -6192
rect 4356 -6210 4365 -6192
rect 4329 -6219 4365 -6210
rect 4563 -6678 4608 -6669
rect 4563 -6696 4572 -6678
rect 4599 -6696 4608 -6678
rect 4626 -6696 4644 -6669
rect 4671 -6696 4680 -6669
rect 4113 -6732 4149 -6723
rect 4113 -6750 4122 -6732
rect 4140 -6750 4149 -6732
rect 4167 -6750 4311 -6723
rect 4329 -6741 4338 -6723
rect 4356 -6741 4365 -6723
rect 4329 -6750 4365 -6741
<< pdiffusion >>
rect 4572 4725 4581 4752
rect 4608 4725 4617 4752
rect 4122 4707 4158 4716
rect 4122 4689 4131 4707
rect 4149 4689 4158 4707
rect 4122 4671 4158 4689
rect 4176 4698 4239 4716
rect 4176 4680 4185 4698
rect 4203 4680 4239 4698
rect 4176 4671 4239 4680
rect 4275 4707 4320 4716
rect 4275 4689 4284 4707
rect 4302 4689 4320 4707
rect 4275 4671 4320 4689
rect 4338 4707 4374 4716
rect 4338 4689 4347 4707
rect 4365 4689 4374 4707
rect 4572 4698 4617 4725
rect 4635 4743 4689 4752
rect 4635 4716 4653 4743
rect 4680 4716 4689 4743
rect 4635 4698 4689 4716
rect 4338 4671 4374 4689
rect 4572 4230 4581 4257
rect 4608 4230 4617 4257
rect 4122 4212 4158 4221
rect 4122 4194 4131 4212
rect 4149 4194 4158 4212
rect 4122 4176 4158 4194
rect 4176 4203 4239 4221
rect 4176 4185 4185 4203
rect 4203 4185 4239 4203
rect 4176 4176 4239 4185
rect 4275 4212 4320 4221
rect 4275 4194 4284 4212
rect 4302 4194 4320 4212
rect 4275 4176 4320 4194
rect 4338 4212 4374 4221
rect 4338 4194 4347 4212
rect 4365 4194 4374 4212
rect 4572 4203 4617 4230
rect 4635 4248 4689 4257
rect 4635 4221 4653 4248
rect 4680 4221 4689 4248
rect 4635 4203 4689 4221
rect 4338 4176 4374 4194
rect 3546 3960 3591 3969
rect 3546 3942 3555 3960
rect 3573 3942 3591 3960
rect 3546 3924 3591 3942
rect 3609 3924 3681 3969
rect 3699 3951 3726 3969
rect 3699 3933 3708 3951
rect 3699 3924 3726 3933
rect 3771 3960 3807 3969
rect 3771 3942 3780 3960
rect 3798 3942 3807 3960
rect 3771 3924 3807 3942
rect 3825 3951 3861 3969
rect 3825 3933 3834 3951
rect 3852 3933 3861 3951
rect 3825 3924 3861 3933
rect 2619 1602 2628 1629
rect 2655 1602 2664 1629
rect 2169 1584 2205 1593
rect 2169 1566 2178 1584
rect 2196 1566 2205 1584
rect 2169 1548 2205 1566
rect 2223 1575 2286 1593
rect 2223 1557 2232 1575
rect 2250 1557 2286 1575
rect 2223 1548 2286 1557
rect 2322 1584 2367 1593
rect 2322 1566 2331 1584
rect 2349 1566 2367 1584
rect 2322 1548 2367 1566
rect 2385 1584 2421 1593
rect 2385 1566 2394 1584
rect 2412 1566 2421 1584
rect 2619 1575 2664 1602
rect 2682 1620 2736 1629
rect 2682 1593 2700 1620
rect 2727 1593 2736 1620
rect 2682 1575 2736 1593
rect 2385 1548 2421 1566
rect 4572 3816 4581 3843
rect 4608 3816 4617 3843
rect 4122 3798 4158 3807
rect 4122 3780 4131 3798
rect 4149 3780 4158 3798
rect 4122 3762 4158 3780
rect 4176 3789 4239 3807
rect 4176 3771 4185 3789
rect 4203 3771 4239 3789
rect 4176 3762 4239 3771
rect 4275 3798 4320 3807
rect 4275 3780 4284 3798
rect 4302 3780 4320 3798
rect 4275 3762 4320 3780
rect 4338 3798 4374 3807
rect 4338 3780 4347 3798
rect 4365 3780 4374 3798
rect 4572 3789 4617 3816
rect 4635 3834 4689 3843
rect 4635 3807 4653 3834
rect 4680 3807 4689 3834
rect 4635 3789 4689 3807
rect 4338 3762 4374 3780
rect 2619 1134 2628 1161
rect 2655 1134 2664 1161
rect 2169 1116 2205 1125
rect 2169 1098 2178 1116
rect 2196 1098 2205 1116
rect 2169 1080 2205 1098
rect 2223 1107 2286 1125
rect 2223 1089 2232 1107
rect 2250 1089 2286 1107
rect 2223 1080 2286 1089
rect 2322 1116 2367 1125
rect 2322 1098 2331 1116
rect 2349 1098 2367 1116
rect 2322 1080 2367 1098
rect 2385 1116 2421 1125
rect 2385 1098 2394 1116
rect 2412 1098 2421 1116
rect 2619 1107 2664 1134
rect 2682 1152 2736 1161
rect 2682 1125 2700 1152
rect 2727 1125 2736 1152
rect 2682 1107 2736 1125
rect 2385 1080 2421 1098
rect 4572 3285 4581 3312
rect 4608 3285 4617 3312
rect 4122 3267 4158 3276
rect 4122 3249 4131 3267
rect 4149 3249 4158 3267
rect 4122 3231 4158 3249
rect 4176 3258 4239 3276
rect 4176 3240 4185 3258
rect 4203 3240 4239 3258
rect 4176 3231 4239 3240
rect 4275 3267 4320 3276
rect 4275 3249 4284 3267
rect 4302 3249 4320 3267
rect 4275 3231 4320 3249
rect 4338 3267 4374 3276
rect 4338 3249 4347 3267
rect 4365 3249 4374 3267
rect 4572 3258 4617 3285
rect 4635 3303 4689 3312
rect 4635 3276 4653 3303
rect 4680 3276 4689 3303
rect 4635 3258 4689 3276
rect 4338 3231 4374 3249
rect 4572 2718 4581 2745
rect 4608 2718 4617 2745
rect 4122 2700 4158 2709
rect 4122 2682 4131 2700
rect 4149 2682 4158 2700
rect 4122 2664 4158 2682
rect 4176 2691 4239 2709
rect 4176 2673 4185 2691
rect 4203 2673 4239 2691
rect 4176 2664 4239 2673
rect 4275 2700 4320 2709
rect 4275 2682 4284 2700
rect 4302 2682 4320 2700
rect 4275 2664 4320 2682
rect 4338 2700 4374 2709
rect 4338 2682 4347 2700
rect 4365 2682 4374 2700
rect 4572 2691 4617 2718
rect 4635 2736 4689 2745
rect 4635 2709 4653 2736
rect 4680 2709 4689 2736
rect 4635 2691 4689 2709
rect 4338 2664 4374 2682
rect 4572 2223 4581 2250
rect 4608 2223 4617 2250
rect 4122 2205 4158 2214
rect 4122 2187 4131 2205
rect 4149 2187 4158 2205
rect 4122 2169 4158 2187
rect 4176 2196 4239 2214
rect 4176 2178 4185 2196
rect 4203 2178 4239 2196
rect 4176 2169 4239 2178
rect 4275 2205 4320 2214
rect 4275 2187 4284 2205
rect 4302 2187 4320 2205
rect 4275 2169 4320 2187
rect 4338 2205 4374 2214
rect 4338 2187 4347 2205
rect 4365 2187 4374 2205
rect 4572 2196 4617 2223
rect 4635 2241 4689 2250
rect 4635 2214 4653 2241
rect 4680 2214 4689 2241
rect 4635 2196 4689 2214
rect 4338 2169 4374 2187
rect 4572 1809 4581 1836
rect 4608 1809 4617 1836
rect 4122 1791 4158 1800
rect 4122 1773 4131 1791
rect 4149 1773 4158 1791
rect 4122 1755 4158 1773
rect 4176 1782 4239 1800
rect 4176 1764 4185 1782
rect 4203 1764 4239 1782
rect 4176 1755 4239 1764
rect 4275 1791 4320 1800
rect 4275 1773 4284 1791
rect 4302 1773 4320 1791
rect 4275 1755 4320 1773
rect 4338 1791 4374 1800
rect 4338 1773 4347 1791
rect 4365 1773 4374 1791
rect 4572 1782 4617 1809
rect 4635 1827 4689 1836
rect 4635 1800 4653 1827
rect 4680 1800 4689 1827
rect 4635 1782 4689 1800
rect 4338 1755 4374 1773
rect 4572 1278 4581 1305
rect 4608 1278 4617 1305
rect 4122 1260 4158 1269
rect 4122 1242 4131 1260
rect 4149 1242 4158 1260
rect 4122 1224 4158 1242
rect 4176 1251 4239 1269
rect 4176 1233 4185 1251
rect 4203 1233 4239 1251
rect 4176 1224 4239 1233
rect 4275 1260 4320 1269
rect 4275 1242 4284 1260
rect 4302 1242 4320 1260
rect 4275 1224 4320 1242
rect 4338 1260 4374 1269
rect 4338 1242 4347 1260
rect 4365 1242 4374 1260
rect 4572 1251 4617 1278
rect 4635 1296 4689 1305
rect 4635 1269 4653 1296
rect 4680 1269 4689 1296
rect 4635 1251 4689 1269
rect 4338 1224 4374 1242
rect 1827 945 1836 972
rect 1863 945 1872 972
rect 1827 918 1872 945
rect 1890 963 1944 972
rect 1890 936 1908 963
rect 1935 936 1944 963
rect 1890 918 1944 936
rect 4563 729 4572 756
rect 4599 729 4608 756
rect 2619 693 2628 720
rect 2655 693 2664 720
rect 2169 675 2205 684
rect 2169 657 2178 675
rect 2196 657 2205 675
rect 1836 621 1845 648
rect 1872 621 1881 648
rect 1836 594 1881 621
rect 1899 639 1953 648
rect 2169 639 2205 657
rect 2223 666 2286 684
rect 2223 648 2232 666
rect 2250 648 2286 666
rect 2223 639 2286 648
rect 2322 675 2367 684
rect 2322 657 2331 675
rect 2349 657 2367 675
rect 2322 639 2367 657
rect 2385 675 2421 684
rect 2385 657 2394 675
rect 2412 657 2421 675
rect 2619 666 2664 693
rect 2682 711 2736 720
rect 2682 684 2700 711
rect 2727 684 2736 711
rect 2682 666 2736 684
rect 4113 711 4149 720
rect 4113 693 4122 711
rect 4140 693 4149 711
rect 4113 675 4149 693
rect 4167 702 4230 720
rect 4167 684 4176 702
rect 4194 684 4230 702
rect 4167 675 4230 684
rect 4266 711 4311 720
rect 4266 693 4275 711
rect 4293 693 4311 711
rect 4266 675 4311 693
rect 4329 711 4365 720
rect 4329 693 4338 711
rect 4356 693 4365 711
rect 4563 702 4608 729
rect 4626 747 4680 756
rect 4626 720 4644 747
rect 4671 720 4680 747
rect 4626 702 4680 720
rect 4329 675 4365 693
rect 2385 639 2421 657
rect 1899 612 1917 639
rect 1944 612 1953 639
rect 1899 594 1953 612
rect 2619 279 2628 306
rect 2655 279 2664 306
rect 2169 261 2205 270
rect 2169 243 2178 261
rect 2196 243 2205 261
rect 2169 225 2205 243
rect 2223 252 2286 270
rect 2223 234 2232 252
rect 2250 234 2286 252
rect 2223 225 2286 234
rect 2322 261 2367 270
rect 2322 243 2331 261
rect 2349 243 2367 261
rect 2322 225 2367 243
rect 2385 261 2421 270
rect 2385 243 2394 261
rect 2412 243 2421 261
rect 2619 252 2664 279
rect 2682 297 2736 306
rect 2682 270 2700 297
rect 2727 270 2736 297
rect 2682 252 2736 270
rect 2385 225 2421 243
rect 4563 234 4572 261
rect 4599 234 4608 261
rect 4113 216 4149 225
rect 4113 198 4122 216
rect 4140 198 4149 216
rect 4113 180 4149 198
rect 4167 207 4230 225
rect 4167 189 4176 207
rect 4194 189 4230 207
rect 4167 180 4230 189
rect 4266 216 4311 225
rect 4266 198 4275 216
rect 4293 198 4311 216
rect 4266 180 4311 198
rect 4329 216 4365 225
rect 4329 198 4338 216
rect 4356 198 4365 216
rect 4563 207 4608 234
rect 4626 252 4680 261
rect 4626 225 4644 252
rect 4671 225 4680 252
rect 4626 207 4680 225
rect 4329 180 4365 198
rect 4563 -180 4572 -153
rect 4599 -180 4608 -153
rect 4113 -198 4149 -189
rect 4113 -216 4122 -198
rect 4140 -216 4149 -198
rect 4113 -234 4149 -216
rect 4167 -207 4230 -189
rect 4167 -225 4176 -207
rect 4194 -225 4230 -207
rect 4167 -234 4230 -225
rect 4266 -198 4311 -189
rect 4266 -216 4275 -198
rect 4293 -216 4311 -198
rect 4266 -234 4311 -216
rect 4329 -198 4365 -189
rect 4329 -216 4338 -198
rect 4356 -216 4365 -198
rect 4563 -207 4608 -180
rect 4626 -162 4680 -153
rect 4626 -189 4644 -162
rect 4671 -189 4680 -162
rect 4626 -207 4680 -189
rect 4329 -234 4365 -216
rect 4563 -711 4572 -684
rect 4599 -711 4608 -684
rect 4113 -729 4149 -720
rect 4113 -747 4122 -729
rect 4140 -747 4149 -729
rect 4113 -765 4149 -747
rect 4167 -738 4230 -720
rect 4167 -756 4176 -738
rect 4194 -756 4230 -738
rect 4167 -765 4230 -756
rect 4266 -729 4311 -720
rect 4266 -747 4275 -729
rect 4293 -747 4311 -729
rect 4266 -765 4311 -747
rect 4329 -729 4365 -720
rect 4329 -747 4338 -729
rect 4356 -747 4365 -729
rect 4563 -738 4608 -711
rect 4626 -693 4680 -684
rect 4626 -720 4644 -693
rect 4671 -720 4680 -693
rect 4626 -738 4680 -720
rect 4329 -765 4365 -747
rect 4563 -1188 4572 -1161
rect 4599 -1188 4608 -1161
rect 4113 -1206 4149 -1197
rect 4113 -1224 4122 -1206
rect 4140 -1224 4149 -1206
rect 4113 -1242 4149 -1224
rect 4167 -1215 4230 -1197
rect 4167 -1233 4176 -1215
rect 4194 -1233 4230 -1215
rect 4167 -1242 4230 -1233
rect 4266 -1206 4311 -1197
rect 4266 -1224 4275 -1206
rect 4293 -1224 4311 -1206
rect 4266 -1242 4311 -1224
rect 4329 -1206 4365 -1197
rect 4329 -1224 4338 -1206
rect 4356 -1224 4365 -1206
rect 4563 -1215 4608 -1188
rect 4626 -1170 4680 -1161
rect 4626 -1197 4644 -1170
rect 4671 -1197 4680 -1170
rect 4626 -1215 4680 -1197
rect 4329 -1242 4365 -1224
rect 4563 -1683 4572 -1656
rect 4599 -1683 4608 -1656
rect 4113 -1701 4149 -1692
rect 4113 -1719 4122 -1701
rect 4140 -1719 4149 -1701
rect 4113 -1737 4149 -1719
rect 4167 -1710 4230 -1692
rect 4167 -1728 4176 -1710
rect 4194 -1728 4230 -1710
rect 4167 -1737 4230 -1728
rect 4266 -1701 4311 -1692
rect 4266 -1719 4275 -1701
rect 4293 -1719 4311 -1701
rect 4266 -1737 4311 -1719
rect 4329 -1701 4365 -1692
rect 4329 -1719 4338 -1701
rect 4356 -1719 4365 -1701
rect 4563 -1710 4608 -1683
rect 4626 -1665 4680 -1656
rect 4626 -1692 4644 -1665
rect 4671 -1692 4680 -1665
rect 4626 -1710 4680 -1692
rect 4329 -1737 4365 -1719
rect 4563 -2097 4572 -2070
rect 4599 -2097 4608 -2070
rect 4113 -2115 4149 -2106
rect 4113 -2133 4122 -2115
rect 4140 -2133 4149 -2115
rect 4113 -2151 4149 -2133
rect 4167 -2124 4230 -2106
rect 4167 -2142 4176 -2124
rect 4194 -2142 4230 -2124
rect 4167 -2151 4230 -2142
rect 4266 -2115 4311 -2106
rect 4266 -2133 4275 -2115
rect 4293 -2133 4311 -2115
rect 4266 -2151 4311 -2133
rect 4329 -2115 4365 -2106
rect 4329 -2133 4338 -2115
rect 4356 -2133 4365 -2115
rect 4563 -2124 4608 -2097
rect 4626 -2079 4680 -2070
rect 4626 -2106 4644 -2079
rect 4671 -2106 4680 -2079
rect 4626 -2124 4680 -2106
rect 4329 -2151 4365 -2133
rect 4563 -2628 4572 -2601
rect 4599 -2628 4608 -2601
rect 4113 -2646 4149 -2637
rect 4113 -2664 4122 -2646
rect 4140 -2664 4149 -2646
rect 4113 -2682 4149 -2664
rect 4167 -2655 4230 -2637
rect 4167 -2673 4176 -2655
rect 4194 -2673 4230 -2655
rect 4167 -2682 4230 -2673
rect 4266 -2646 4311 -2637
rect 4266 -2664 4275 -2646
rect 4293 -2664 4311 -2646
rect 4266 -2682 4311 -2664
rect 4329 -2646 4365 -2637
rect 4329 -2664 4338 -2646
rect 4356 -2664 4365 -2646
rect 4563 -2655 4608 -2628
rect 4626 -2610 4680 -2601
rect 4626 -2637 4644 -2610
rect 4671 -2637 4680 -2610
rect 4626 -2655 4680 -2637
rect 4329 -2682 4365 -2664
rect 4563 -3195 4572 -3168
rect 4599 -3195 4608 -3168
rect 4113 -3213 4149 -3204
rect 4113 -3231 4122 -3213
rect 4140 -3231 4149 -3213
rect 4113 -3249 4149 -3231
rect 4167 -3222 4230 -3204
rect 4167 -3240 4176 -3222
rect 4194 -3240 4230 -3222
rect 4167 -3249 4230 -3240
rect 4266 -3213 4311 -3204
rect 4266 -3231 4275 -3213
rect 4293 -3231 4311 -3213
rect 4266 -3249 4311 -3231
rect 4329 -3213 4365 -3204
rect 4329 -3231 4338 -3213
rect 4356 -3231 4365 -3213
rect 4563 -3222 4608 -3195
rect 4626 -3177 4680 -3168
rect 4626 -3204 4644 -3177
rect 4671 -3204 4680 -3177
rect 4626 -3222 4680 -3204
rect 4329 -3249 4365 -3231
rect 4563 -3690 4572 -3663
rect 4599 -3690 4608 -3663
rect 4113 -3708 4149 -3699
rect 4113 -3726 4122 -3708
rect 4140 -3726 4149 -3708
rect 4113 -3744 4149 -3726
rect 4167 -3717 4230 -3699
rect 4167 -3735 4176 -3717
rect 4194 -3735 4230 -3717
rect 4167 -3744 4230 -3735
rect 4266 -3708 4311 -3699
rect 4266 -3726 4275 -3708
rect 4293 -3726 4311 -3708
rect 4266 -3744 4311 -3726
rect 4329 -3708 4365 -3699
rect 4329 -3726 4338 -3708
rect 4356 -3726 4365 -3708
rect 4563 -3717 4608 -3690
rect 4626 -3672 4680 -3663
rect 4626 -3699 4644 -3672
rect 4671 -3699 4680 -3672
rect 4626 -3717 4680 -3699
rect 4329 -3744 4365 -3726
rect 4563 -4104 4572 -4077
rect 4599 -4104 4608 -4077
rect 4113 -4122 4149 -4113
rect 4113 -4140 4122 -4122
rect 4140 -4140 4149 -4122
rect 4113 -4158 4149 -4140
rect 4167 -4131 4230 -4113
rect 4167 -4149 4176 -4131
rect 4194 -4149 4230 -4131
rect 4167 -4158 4230 -4149
rect 4266 -4122 4311 -4113
rect 4266 -4140 4275 -4122
rect 4293 -4140 4311 -4122
rect 4266 -4158 4311 -4140
rect 4329 -4122 4365 -4113
rect 4329 -4140 4338 -4122
rect 4356 -4140 4365 -4122
rect 4563 -4131 4608 -4104
rect 4626 -4086 4680 -4077
rect 4626 -4113 4644 -4086
rect 4671 -4113 4680 -4086
rect 4626 -4131 4680 -4113
rect 4329 -4158 4365 -4140
rect 4563 -4635 4572 -4608
rect 4599 -4635 4608 -4608
rect 4113 -4653 4149 -4644
rect 4113 -4671 4122 -4653
rect 4140 -4671 4149 -4653
rect 4113 -4689 4149 -4671
rect 4167 -4662 4230 -4644
rect 4167 -4680 4176 -4662
rect 4194 -4680 4230 -4662
rect 4167 -4689 4230 -4680
rect 4266 -4653 4311 -4644
rect 4266 -4671 4275 -4653
rect 4293 -4671 4311 -4653
rect 4266 -4689 4311 -4671
rect 4329 -4653 4365 -4644
rect 4329 -4671 4338 -4653
rect 4356 -4671 4365 -4653
rect 4563 -4662 4608 -4635
rect 4626 -4617 4680 -4608
rect 4626 -4644 4644 -4617
rect 4671 -4644 4680 -4617
rect 4626 -4662 4680 -4644
rect 4329 -4689 4365 -4671
rect 4563 -5130 4572 -5103
rect 4599 -5130 4608 -5103
rect 4113 -5148 4149 -5139
rect 4113 -5166 4122 -5148
rect 4140 -5166 4149 -5148
rect 4113 -5184 4149 -5166
rect 4167 -5157 4230 -5139
rect 4167 -5175 4176 -5157
rect 4194 -5175 4230 -5157
rect 4167 -5184 4230 -5175
rect 4266 -5148 4311 -5139
rect 4266 -5166 4275 -5148
rect 4293 -5166 4311 -5148
rect 4266 -5184 4311 -5166
rect 4329 -5148 4365 -5139
rect 4329 -5166 4338 -5148
rect 4356 -5166 4365 -5148
rect 4563 -5157 4608 -5130
rect 4626 -5112 4680 -5103
rect 4626 -5139 4644 -5112
rect 4671 -5139 4680 -5112
rect 4626 -5157 4680 -5139
rect 4329 -5184 4365 -5166
rect 4563 -5625 4572 -5598
rect 4599 -5625 4608 -5598
rect 4113 -5643 4149 -5634
rect 4113 -5661 4122 -5643
rect 4140 -5661 4149 -5643
rect 4113 -5679 4149 -5661
rect 4167 -5652 4230 -5634
rect 4167 -5670 4176 -5652
rect 4194 -5670 4230 -5652
rect 4167 -5679 4230 -5670
rect 4266 -5643 4311 -5634
rect 4266 -5661 4275 -5643
rect 4293 -5661 4311 -5643
rect 4266 -5679 4311 -5661
rect 4329 -5643 4365 -5634
rect 4329 -5661 4338 -5643
rect 4356 -5661 4365 -5643
rect 4563 -5652 4608 -5625
rect 4626 -5607 4680 -5598
rect 4626 -5634 4644 -5607
rect 4671 -5634 4680 -5607
rect 4626 -5652 4680 -5634
rect 4329 -5679 4365 -5661
rect 4563 -6039 4572 -6012
rect 4599 -6039 4608 -6012
rect 4113 -6057 4149 -6048
rect 4113 -6075 4122 -6057
rect 4140 -6075 4149 -6057
rect 4113 -6093 4149 -6075
rect 4167 -6066 4230 -6048
rect 4167 -6084 4176 -6066
rect 4194 -6084 4230 -6066
rect 4167 -6093 4230 -6084
rect 4266 -6057 4311 -6048
rect 4266 -6075 4275 -6057
rect 4293 -6075 4311 -6057
rect 4266 -6093 4311 -6075
rect 4329 -6057 4365 -6048
rect 4329 -6075 4338 -6057
rect 4356 -6075 4365 -6057
rect 4563 -6066 4608 -6039
rect 4626 -6021 4680 -6012
rect 4626 -6048 4644 -6021
rect 4671 -6048 4680 -6021
rect 4626 -6066 4680 -6048
rect 4329 -6093 4365 -6075
rect 4563 -6570 4572 -6543
rect 4599 -6570 4608 -6543
rect 4113 -6588 4149 -6579
rect 4113 -6606 4122 -6588
rect 4140 -6606 4149 -6588
rect 4113 -6624 4149 -6606
rect 4167 -6597 4230 -6579
rect 4167 -6615 4176 -6597
rect 4194 -6615 4230 -6597
rect 4167 -6624 4230 -6615
rect 4266 -6588 4311 -6579
rect 4266 -6606 4275 -6588
rect 4293 -6606 4311 -6588
rect 4266 -6624 4311 -6606
rect 4329 -6588 4365 -6579
rect 4329 -6606 4338 -6588
rect 4356 -6606 4365 -6588
rect 4563 -6597 4608 -6570
rect 4626 -6552 4680 -6543
rect 4626 -6579 4644 -6552
rect 4671 -6579 4680 -6552
rect 4626 -6597 4680 -6579
rect 4329 -6624 4365 -6606
<< ndcontact >>
rect 4581 4590 4608 4617
rect 4653 4599 4680 4626
rect 4131 4545 4149 4563
rect 4347 4554 4365 4572
rect 4581 4095 4608 4122
rect 4653 4104 4680 4131
rect 4131 4050 4149 4068
rect 4347 4059 4365 4077
rect 3564 3816 3582 3834
rect 3618 3816 3636 3834
rect 3654 3816 3672 3834
rect 3708 3816 3726 3834
rect 3780 3816 3798 3834
rect 3834 3816 3852 3834
rect 2628 1467 2655 1494
rect 2700 1476 2727 1503
rect 2178 1422 2196 1440
rect 2394 1431 2412 1449
rect 4581 3681 4608 3708
rect 4653 3690 4680 3717
rect 4131 3636 4149 3654
rect 4347 3645 4365 3663
rect 4581 3150 4608 3177
rect 4653 3159 4680 3186
rect 4131 3105 4149 3123
rect 4347 3114 4365 3132
rect 4581 2583 4608 2610
rect 4653 2592 4680 2619
rect 4131 2538 4149 2556
rect 4347 2547 4365 2565
rect 4581 2088 4608 2115
rect 4653 2097 4680 2124
rect 4131 2043 4149 2061
rect 4347 2052 4365 2070
rect 4581 1674 4608 1701
rect 4653 1683 4680 1710
rect 4131 1629 4149 1647
rect 4347 1638 4365 1656
rect 4581 1143 4608 1170
rect 4653 1152 4680 1179
rect 4131 1098 4149 1116
rect 4347 1107 4365 1125
rect 2628 999 2655 1026
rect 2700 1008 2727 1035
rect 2178 954 2196 972
rect 2394 963 2412 981
rect 1836 810 1863 837
rect 1908 819 1935 846
rect 2628 558 2655 585
rect 2700 567 2727 594
rect 1845 486 1872 513
rect 1917 495 1944 522
rect 2178 513 2196 531
rect 2394 522 2412 540
rect 2628 144 2655 171
rect 2700 153 2727 180
rect 2178 99 2196 117
rect 2394 108 2412 126
rect 4572 594 4599 621
rect 4644 603 4671 630
rect 4122 549 4140 567
rect 4338 558 4356 576
rect 4572 99 4599 126
rect 4644 108 4671 135
rect 4122 54 4140 72
rect 4338 63 4356 81
rect 4572 -315 4599 -288
rect 4644 -306 4671 -279
rect 4122 -360 4140 -342
rect 4338 -351 4356 -333
rect 4572 -846 4599 -819
rect 4644 -837 4671 -810
rect 4122 -891 4140 -873
rect 4338 -882 4356 -864
rect 4572 -1323 4599 -1296
rect 4644 -1314 4671 -1287
rect 4122 -1368 4140 -1350
rect 4338 -1359 4356 -1341
rect 4572 -1818 4599 -1791
rect 4644 -1809 4671 -1782
rect 4122 -1863 4140 -1845
rect 4338 -1854 4356 -1836
rect 4572 -2232 4599 -2205
rect 4644 -2223 4671 -2196
rect 4122 -2277 4140 -2259
rect 4338 -2268 4356 -2250
rect 4572 -2763 4599 -2736
rect 4644 -2754 4671 -2727
rect 4122 -2808 4140 -2790
rect 4338 -2799 4356 -2781
rect 4572 -3330 4599 -3303
rect 4644 -3321 4671 -3294
rect 4122 -3375 4140 -3357
rect 4338 -3366 4356 -3348
rect 4572 -3825 4599 -3798
rect 4644 -3816 4671 -3789
rect 4122 -3870 4140 -3852
rect 4338 -3861 4356 -3843
rect 4572 -4239 4599 -4212
rect 4644 -4230 4671 -4203
rect 4122 -4284 4140 -4266
rect 4338 -4275 4356 -4257
rect 4572 -4770 4599 -4743
rect 4644 -4761 4671 -4734
rect 4122 -4815 4140 -4797
rect 4338 -4806 4356 -4788
rect 4572 -5265 4599 -5238
rect 4644 -5256 4671 -5229
rect 4122 -5310 4140 -5292
rect 4338 -5301 4356 -5283
rect 4572 -5760 4599 -5733
rect 4644 -5751 4671 -5724
rect 4122 -5805 4140 -5787
rect 4338 -5796 4356 -5778
rect 4572 -6174 4599 -6147
rect 4644 -6165 4671 -6138
rect 4122 -6219 4140 -6201
rect 4338 -6210 4356 -6192
rect 4572 -6705 4599 -6678
rect 4644 -6696 4671 -6669
rect 4122 -6750 4140 -6732
rect 4338 -6741 4356 -6723
<< pdcontact >>
rect 4581 4725 4608 4752
rect 4131 4689 4149 4707
rect 4185 4680 4203 4698
rect 4284 4689 4302 4707
rect 4347 4689 4365 4707
rect 4653 4716 4680 4743
rect 4581 4230 4608 4257
rect 4131 4194 4149 4212
rect 4185 4185 4203 4203
rect 4284 4194 4302 4212
rect 4347 4194 4365 4212
rect 4653 4221 4680 4248
rect 3555 3942 3573 3960
rect 3708 3933 3726 3951
rect 3780 3942 3798 3960
rect 3834 3933 3852 3951
rect 2628 1602 2655 1629
rect 2178 1566 2196 1584
rect 2232 1557 2250 1575
rect 2331 1566 2349 1584
rect 2394 1566 2412 1584
rect 2700 1593 2727 1620
rect 4581 3816 4608 3843
rect 4131 3780 4149 3798
rect 4185 3771 4203 3789
rect 4284 3780 4302 3798
rect 4347 3780 4365 3798
rect 4653 3807 4680 3834
rect 2628 1134 2655 1161
rect 2178 1098 2196 1116
rect 2232 1089 2250 1107
rect 2331 1098 2349 1116
rect 2394 1098 2412 1116
rect 2700 1125 2727 1152
rect 4581 3285 4608 3312
rect 4131 3249 4149 3267
rect 4185 3240 4203 3258
rect 4284 3249 4302 3267
rect 4347 3249 4365 3267
rect 4653 3276 4680 3303
rect 4581 2718 4608 2745
rect 4131 2682 4149 2700
rect 4185 2673 4203 2691
rect 4284 2682 4302 2700
rect 4347 2682 4365 2700
rect 4653 2709 4680 2736
rect 4581 2223 4608 2250
rect 4131 2187 4149 2205
rect 4185 2178 4203 2196
rect 4284 2187 4302 2205
rect 4347 2187 4365 2205
rect 4653 2214 4680 2241
rect 4581 1809 4608 1836
rect 4131 1773 4149 1791
rect 4185 1764 4203 1782
rect 4284 1773 4302 1791
rect 4347 1773 4365 1791
rect 4653 1800 4680 1827
rect 4581 1278 4608 1305
rect 4131 1242 4149 1260
rect 4185 1233 4203 1251
rect 4284 1242 4302 1260
rect 4347 1242 4365 1260
rect 4653 1269 4680 1296
rect 1836 945 1863 972
rect 1908 936 1935 963
rect 4572 729 4599 756
rect 2628 693 2655 720
rect 2178 657 2196 675
rect 1845 621 1872 648
rect 2232 648 2250 666
rect 2331 657 2349 675
rect 2394 657 2412 675
rect 2700 684 2727 711
rect 4122 693 4140 711
rect 4176 684 4194 702
rect 4275 693 4293 711
rect 4338 693 4356 711
rect 4644 720 4671 747
rect 1917 612 1944 639
rect 2628 279 2655 306
rect 2178 243 2196 261
rect 2232 234 2250 252
rect 2331 243 2349 261
rect 2394 243 2412 261
rect 2700 270 2727 297
rect 4572 234 4599 261
rect 4122 198 4140 216
rect 4176 189 4194 207
rect 4275 198 4293 216
rect 4338 198 4356 216
rect 4644 225 4671 252
rect 4572 -180 4599 -153
rect 4122 -216 4140 -198
rect 4176 -225 4194 -207
rect 4275 -216 4293 -198
rect 4338 -216 4356 -198
rect 4644 -189 4671 -162
rect 4572 -711 4599 -684
rect 4122 -747 4140 -729
rect 4176 -756 4194 -738
rect 4275 -747 4293 -729
rect 4338 -747 4356 -729
rect 4644 -720 4671 -693
rect 4572 -1188 4599 -1161
rect 4122 -1224 4140 -1206
rect 4176 -1233 4194 -1215
rect 4275 -1224 4293 -1206
rect 4338 -1224 4356 -1206
rect 4644 -1197 4671 -1170
rect 4572 -1683 4599 -1656
rect 4122 -1719 4140 -1701
rect 4176 -1728 4194 -1710
rect 4275 -1719 4293 -1701
rect 4338 -1719 4356 -1701
rect 4644 -1692 4671 -1665
rect 4572 -2097 4599 -2070
rect 4122 -2133 4140 -2115
rect 4176 -2142 4194 -2124
rect 4275 -2133 4293 -2115
rect 4338 -2133 4356 -2115
rect 4644 -2106 4671 -2079
rect 4572 -2628 4599 -2601
rect 4122 -2664 4140 -2646
rect 4176 -2673 4194 -2655
rect 4275 -2664 4293 -2646
rect 4338 -2664 4356 -2646
rect 4644 -2637 4671 -2610
rect 4572 -3195 4599 -3168
rect 4122 -3231 4140 -3213
rect 4176 -3240 4194 -3222
rect 4275 -3231 4293 -3213
rect 4338 -3231 4356 -3213
rect 4644 -3204 4671 -3177
rect 4572 -3690 4599 -3663
rect 4122 -3726 4140 -3708
rect 4176 -3735 4194 -3717
rect 4275 -3726 4293 -3708
rect 4338 -3726 4356 -3708
rect 4644 -3699 4671 -3672
rect 4572 -4104 4599 -4077
rect 4122 -4140 4140 -4122
rect 4176 -4149 4194 -4131
rect 4275 -4140 4293 -4122
rect 4338 -4140 4356 -4122
rect 4644 -4113 4671 -4086
rect 4572 -4635 4599 -4608
rect 4122 -4671 4140 -4653
rect 4176 -4680 4194 -4662
rect 4275 -4671 4293 -4653
rect 4338 -4671 4356 -4653
rect 4644 -4644 4671 -4617
rect 4572 -5130 4599 -5103
rect 4122 -5166 4140 -5148
rect 4176 -5175 4194 -5157
rect 4275 -5166 4293 -5148
rect 4338 -5166 4356 -5148
rect 4644 -5139 4671 -5112
rect 4572 -5625 4599 -5598
rect 4122 -5661 4140 -5643
rect 4176 -5670 4194 -5652
rect 4275 -5661 4293 -5643
rect 4338 -5661 4356 -5643
rect 4644 -5634 4671 -5607
rect 4572 -6039 4599 -6012
rect 4122 -6075 4140 -6057
rect 4176 -6084 4194 -6066
rect 4275 -6075 4293 -6057
rect 4338 -6075 4356 -6057
rect 4644 -6048 4671 -6021
rect 4572 -6570 4599 -6543
rect 4122 -6606 4140 -6588
rect 4176 -6615 4194 -6597
rect 4275 -6606 4293 -6588
rect 4338 -6606 4356 -6588
rect 4644 -6579 4671 -6552
<< polysilicon >>
rect 846 4860 4338 4878
rect 846 -162 864 4860
rect 4158 4716 4176 4743
rect 4320 4716 4338 4860
rect 4617 4752 4635 4869
rect 4158 4608 4176 4671
rect 3987 4590 4176 4608
rect 3987 4113 4005 4590
rect 4158 4572 4176 4590
rect 4320 4572 4338 4671
rect 4617 4662 4635 4698
rect 4626 4635 4635 4662
rect 4617 4626 4635 4635
rect 4617 4581 4635 4599
rect 4158 4536 4176 4545
rect 4320 4536 4338 4545
rect 4158 4221 4176 4248
rect 4320 4221 4338 4356
rect 4617 4257 4635 4374
rect 4158 4113 4176 4176
rect 3987 4095 4176 4113
rect 3591 3969 3609 3987
rect 3681 3969 3699 3987
rect 3807 3969 3825 3987
rect 3591 3861 3609 3924
rect 3015 3843 3609 3861
rect 2664 1629 2682 1746
rect 2205 1593 2223 1620
rect 2367 1593 2385 1620
rect 2205 1494 2223 1548
rect 2367 1476 2385 1548
rect 2664 1539 2682 1575
rect 3015 1548 3033 3843
rect 3591 3834 3609 3843
rect 3681 3834 3699 3924
rect 3807 3879 3825 3924
rect 3987 3879 4005 4095
rect 4158 4077 4176 4095
rect 4320 4077 4338 4176
rect 4617 4167 4635 4203
rect 4626 4140 4635 4167
rect 4617 4131 4635 4140
rect 4617 4086 4635 4104
rect 4158 4041 4176 4050
rect 4320 4041 4338 4050
rect 3816 3861 3825 3879
rect 3897 3861 4005 3879
rect 3807 3834 3825 3861
rect 3591 3798 3609 3807
rect 3681 3510 3699 3807
rect 3807 3798 3825 3807
rect 2673 1512 2682 1539
rect 2763 1521 3033 1548
rect 3114 3492 3699 3510
rect 3987 3690 4005 3861
rect 4617 3843 4635 3960
rect 4158 3807 4176 3834
rect 4320 3807 4338 3834
rect 4158 3690 4176 3762
rect 3987 3672 4176 3690
rect 2664 1503 2682 1512
rect 2205 1449 2223 1476
rect 2664 1458 2682 1476
rect 2367 1449 2385 1458
rect 2205 1413 2223 1422
rect 2367 1413 2385 1422
rect 1737 1161 2133 1179
rect 2664 1161 2682 1278
rect 1737 882 1755 1161
rect 2115 1017 2133 1161
rect 2205 1125 2223 1152
rect 2367 1125 2385 1152
rect 2205 1017 2223 1080
rect 2115 999 2223 1017
rect 1872 972 1890 990
rect 2205 981 2223 999
rect 2367 1008 2385 1080
rect 2664 1071 2682 1107
rect 3114 1080 3132 3492
rect 3987 3168 4005 3672
rect 4158 3663 4176 3672
rect 4320 3663 4338 3762
rect 4617 3753 4635 3789
rect 4626 3726 4635 3753
rect 4617 3717 4635 3726
rect 4617 3672 4635 3690
rect 4158 3627 4176 3636
rect 4320 3546 4338 3636
rect 4617 3312 4635 3429
rect 4158 3276 4176 3303
rect 4320 3276 4338 3303
rect 4158 3168 4176 3231
rect 3987 3150 4176 3168
rect 3987 2601 4005 3150
rect 4158 3132 4176 3150
rect 4320 3132 4338 3231
rect 4617 3222 4635 3258
rect 4626 3195 4635 3222
rect 4617 3186 4635 3195
rect 4617 3141 4635 3159
rect 4158 3096 4176 3105
rect 4320 3006 4338 3105
rect 4617 2745 4635 2862
rect 4158 2709 4176 2736
rect 4320 2709 4338 2736
rect 4158 2601 4176 2664
rect 3987 2583 4176 2601
rect 3987 2106 4005 2583
rect 4158 2565 4176 2583
rect 4320 2565 4338 2664
rect 4617 2655 4635 2691
rect 4626 2628 4635 2655
rect 4617 2619 4635 2628
rect 4617 2574 4635 2592
rect 4158 2529 4176 2538
rect 4320 2448 4338 2538
rect 4617 2250 4635 2367
rect 4158 2214 4176 2241
rect 4320 2214 4338 2241
rect 4158 2106 4176 2169
rect 3987 2088 4176 2106
rect 3987 1872 4005 2088
rect 4158 2070 4176 2088
rect 4320 2070 4338 2169
rect 4617 2160 4635 2196
rect 4626 2133 4635 2160
rect 4617 2124 4635 2133
rect 4617 2079 4635 2097
rect 4158 2034 4176 2043
rect 4320 1971 4338 2043
rect 3978 1854 4005 1872
rect 3987 1683 4005 1854
rect 4617 1836 4635 1953
rect 4158 1800 4176 1827
rect 4320 1800 4338 1827
rect 4158 1683 4176 1755
rect 3987 1665 4176 1683
rect 3987 1161 4005 1665
rect 4158 1656 4176 1665
rect 4320 1656 4338 1755
rect 4617 1746 4635 1782
rect 4626 1719 4635 1746
rect 4617 1710 4635 1719
rect 4617 1665 4635 1683
rect 4158 1620 4176 1629
rect 4320 1530 4338 1629
rect 4617 1305 4635 1422
rect 4158 1269 4176 1296
rect 4320 1269 4338 1296
rect 4158 1161 4176 1224
rect 3987 1143 4176 1161
rect 4158 1125 4176 1143
rect 4320 1125 4338 1224
rect 4617 1215 4635 1251
rect 4626 1188 4635 1215
rect 4617 1179 4635 1188
rect 4617 1134 4635 1152
rect 4158 1089 4176 1098
rect 2673 1044 2682 1071
rect 2763 1053 3132 1080
rect 2664 1035 2682 1044
rect 4320 1026 4338 1098
rect 2664 990 2682 1008
rect 2367 981 2385 990
rect 2205 945 2223 954
rect 2367 945 2385 954
rect 1872 882 1890 918
rect 1620 855 1890 882
rect 1620 18 1638 855
rect 1872 846 1890 855
rect 1872 801 1890 819
rect 2664 720 2682 837
rect 4608 756 4626 873
rect 4149 720 4167 747
rect 4311 720 4329 747
rect 2205 684 2223 711
rect 2367 684 2385 711
rect 1881 648 1899 666
rect 2205 594 2223 639
rect 1881 558 1899 594
rect 1674 531 1899 558
rect 2205 540 2223 576
rect 2367 567 2385 639
rect 2664 630 2682 666
rect 2673 603 2682 630
rect 2763 612 3996 639
rect 4149 612 4167 675
rect 2664 594 2682 603
rect 3978 594 4167 612
rect 2340 549 2385 567
rect 2664 549 2682 567
rect 2340 540 2358 549
rect 2367 540 2385 549
rect 1674 414 1692 531
rect 1881 522 1899 531
rect 2205 504 2223 513
rect 1881 477 1899 495
rect 2340 414 2358 513
rect 2367 504 2385 513
rect 1674 396 2358 414
rect 2061 189 2079 396
rect 2664 306 2682 423
rect 2205 270 2223 297
rect 2367 270 2385 297
rect 2205 189 2223 225
rect 2061 171 2223 189
rect 2205 126 2223 171
rect 2367 153 2385 225
rect 2664 216 2682 252
rect 2673 189 2682 216
rect 2664 180 2682 189
rect 2322 135 2385 153
rect 2664 135 2682 153
rect 2322 126 2340 135
rect 2367 126 2385 135
rect 2754 99 3087 117
rect 2205 90 2223 99
rect 2322 18 2340 99
rect 2367 90 2385 99
rect 1620 0 2340 18
rect 3069 72 3087 99
rect 3762 -162 3780 450
rect 846 -180 3780 -162
rect 3978 117 3996 594
rect 4149 576 4167 594
rect 4311 576 4329 675
rect 4608 666 4626 702
rect 4617 639 4626 666
rect 4608 630 4626 639
rect 4608 585 4626 603
rect 4149 540 4167 549
rect 4311 468 4329 549
rect 4608 261 4626 378
rect 4149 225 4167 252
rect 4311 225 4329 252
rect 4149 117 4167 180
rect 3978 99 4167 117
rect 846 -3447 864 -180
rect 3978 -306 3996 99
rect 4149 81 4167 99
rect 4311 81 4329 180
rect 4608 171 4626 207
rect 4617 144 4626 171
rect 4608 135 4626 144
rect 4608 90 4626 108
rect 4149 45 4167 54
rect 4311 -27 4329 54
rect 4608 -153 4626 -36
rect 4149 -189 4167 -162
rect 4311 -189 4329 -162
rect 4149 -306 4167 -234
rect 3978 -324 4167 -306
rect 1035 -981 1053 -387
rect 3978 -828 3996 -324
rect 4149 -333 4167 -324
rect 4311 -333 4329 -234
rect 4608 -243 4626 -207
rect 4617 -270 4626 -243
rect 4608 -279 4626 -270
rect 4608 -324 4626 -306
rect 4149 -369 4167 -360
rect 4311 -468 4329 -360
rect 4608 -684 4626 -567
rect 4149 -720 4167 -693
rect 4311 -720 4329 -693
rect 4149 -828 4167 -765
rect 3978 -846 4167 -828
rect 1035 -4509 1053 -1035
rect 3978 -1305 3996 -846
rect 4149 -864 4167 -846
rect 4311 -864 4329 -765
rect 4608 -774 4626 -738
rect 4617 -801 4626 -774
rect 4608 -810 4626 -801
rect 4608 -855 4626 -837
rect 4149 -900 4167 -891
rect 4311 -990 4329 -891
rect 4608 -1161 4626 -1044
rect 4149 -1197 4167 -1170
rect 4311 -1197 4329 -1170
rect 4149 -1305 4167 -1242
rect 3978 -1323 4167 -1305
rect 3978 -1800 3996 -1323
rect 4149 -1341 4167 -1323
rect 4311 -1341 4329 -1242
rect 4608 -1251 4626 -1215
rect 4617 -1278 4626 -1251
rect 4608 -1287 4626 -1278
rect 4608 -1332 4626 -1314
rect 4149 -1377 4167 -1368
rect 4311 -1440 4329 -1368
rect 4608 -1656 4626 -1539
rect 4149 -1692 4167 -1665
rect 4311 -1692 4329 -1665
rect 4149 -1800 4167 -1737
rect 3978 -1818 4167 -1800
rect 3978 -2223 3996 -1818
rect 4149 -1836 4167 -1818
rect 4311 -1836 4329 -1737
rect 4608 -1746 4626 -1710
rect 4617 -1773 4626 -1746
rect 4608 -1782 4626 -1773
rect 4608 -1827 4626 -1809
rect 4149 -1872 4167 -1863
rect 4311 -1935 4329 -1863
rect 4608 -2070 4626 -1953
rect 4149 -2106 4167 -2079
rect 4311 -2106 4329 -2079
rect 4149 -2223 4167 -2151
rect 3978 -2241 4167 -2223
rect 3978 -2745 3996 -2241
rect 4149 -2250 4167 -2241
rect 4311 -2250 4329 -2151
rect 4608 -2160 4626 -2124
rect 4617 -2187 4626 -2160
rect 4608 -2196 4626 -2187
rect 4608 -2241 4626 -2223
rect 4149 -2286 4167 -2277
rect 4311 -2322 4329 -2277
rect 4608 -2601 4626 -2484
rect 4149 -2637 4167 -2610
rect 4311 -2637 4329 -2610
rect 4149 -2745 4167 -2682
rect 3978 -2763 4167 -2745
rect 4149 -2781 4167 -2763
rect 4311 -2781 4329 -2682
rect 4608 -2691 4626 -2655
rect 4617 -2718 4626 -2691
rect 4608 -2727 4626 -2718
rect 4608 -2772 4626 -2754
rect 4149 -2817 4167 -2808
rect 4311 -2889 4329 -2808
rect 4608 -3168 4626 -3051
rect 4149 -3204 4167 -3177
rect 4311 -3204 4329 -3177
rect 4149 -3312 4167 -3249
rect 3978 -3321 4167 -3312
rect 4014 -3330 4167 -3321
rect 4149 -3348 4167 -3330
rect 4311 -3348 4329 -3249
rect 4608 -3258 4626 -3222
rect 4617 -3285 4626 -3258
rect 4608 -3294 4626 -3285
rect 4608 -3339 4626 -3321
rect 3978 -3807 3996 -3348
rect 4149 -3384 4167 -3375
rect 4311 -3447 4329 -3375
rect 4608 -3663 4626 -3546
rect 4149 -3699 4167 -3672
rect 4311 -3699 4329 -3672
rect 4149 -3807 4167 -3744
rect 3978 -3825 4167 -3807
rect 3978 -4230 3996 -3825
rect 4149 -3843 4167 -3825
rect 4311 -3843 4329 -3744
rect 4608 -3753 4626 -3717
rect 4617 -3780 4626 -3753
rect 4608 -3789 4626 -3780
rect 4608 -3834 4626 -3816
rect 4149 -3879 4167 -3870
rect 4311 -3960 4329 -3870
rect 4608 -4077 4626 -3960
rect 4149 -4113 4167 -4086
rect 4311 -4113 4329 -4086
rect 4149 -4230 4167 -4158
rect 3978 -4248 4167 -4230
rect 3978 -4752 3996 -4248
rect 4149 -4257 4167 -4248
rect 4311 -4257 4329 -4158
rect 4608 -4167 4626 -4131
rect 4617 -4194 4626 -4167
rect 4608 -4203 4626 -4194
rect 4608 -4248 4626 -4230
rect 4149 -4293 4167 -4284
rect 4311 -4392 4329 -4284
rect 4608 -4608 4626 -4491
rect 4149 -4644 4167 -4617
rect 4311 -4644 4329 -4617
rect 4149 -4752 4167 -4689
rect 3978 -4770 4167 -4752
rect 3978 -5247 3996 -4770
rect 4149 -4788 4167 -4770
rect 4311 -4788 4329 -4689
rect 4608 -4698 4626 -4662
rect 4617 -4725 4626 -4698
rect 4608 -4734 4626 -4725
rect 4608 -4779 4626 -4761
rect 4149 -4824 4167 -4815
rect 4311 -4905 4329 -4815
rect 4608 -5103 4626 -4986
rect 4149 -5139 4167 -5112
rect 4311 -5139 4329 -5112
rect 4149 -5247 4167 -5184
rect 3978 -5265 4167 -5247
rect 3978 -5742 3996 -5265
rect 4149 -5283 4167 -5265
rect 4311 -5283 4329 -5184
rect 4608 -5193 4626 -5157
rect 4617 -5220 4626 -5193
rect 4608 -5229 4626 -5220
rect 4608 -5274 4626 -5256
rect 4149 -5319 4167 -5310
rect 4311 -5382 4329 -5310
rect 4608 -5598 4626 -5481
rect 4149 -5634 4167 -5607
rect 4311 -5634 4329 -5607
rect 4149 -5742 4167 -5679
rect 3978 -5760 4167 -5742
rect 3978 -6165 3996 -5760
rect 4149 -5778 4167 -5760
rect 4311 -5778 4329 -5679
rect 4608 -5688 4626 -5652
rect 4617 -5715 4626 -5688
rect 4608 -5724 4626 -5715
rect 4608 -5769 4626 -5751
rect 4149 -5814 4167 -5805
rect 4311 -5868 4329 -5805
rect 4608 -6012 4626 -5895
rect 4149 -6048 4167 -6021
rect 4311 -6048 4329 -6021
rect 4149 -6165 4167 -6093
rect 3978 -6183 4167 -6165
rect 3978 -6687 3996 -6183
rect 4149 -6192 4167 -6183
rect 4311 -6192 4329 -6093
rect 4608 -6102 4626 -6066
rect 4617 -6129 4626 -6102
rect 4608 -6138 4626 -6129
rect 4608 -6183 4626 -6165
rect 4149 -6228 4167 -6219
rect 4311 -6300 4329 -6219
rect 4608 -6543 4626 -6426
rect 4149 -6579 4167 -6552
rect 4311 -6579 4329 -6552
rect 4149 -6687 4167 -6624
rect 3978 -6705 4167 -6687
rect 4149 -6723 4167 -6705
rect 4311 -6723 4329 -6624
rect 4608 -6633 4626 -6597
rect 4617 -6660 4626 -6633
rect 4608 -6669 4626 -6660
rect 4608 -6714 4626 -6696
rect 4149 -6759 4167 -6750
rect 4311 -6822 4329 -6750
rect 3591 -6840 4329 -6822
<< polycontact >>
rect 4599 4635 4626 4662
rect 4320 4356 4338 4374
rect 2196 1476 2223 1494
rect 4599 4140 4626 4167
rect 3807 3861 3816 3879
rect 3852 3861 3897 3879
rect 2646 1512 2673 1539
rect 2727 1521 2763 1548
rect 2349 1458 2385 1476
rect 4599 3726 4626 3753
rect 4320 3528 4338 3546
rect 4599 3195 4626 3222
rect 4320 2988 4338 3006
rect 4599 2628 4626 2655
rect 4311 2412 4347 2448
rect 4599 2133 4626 2160
rect 4311 1935 4347 1971
rect 4599 1719 4626 1746
rect 4302 1494 4347 1530
rect 4599 1188 4626 1215
rect 2646 1044 2673 1071
rect 2718 1053 2763 1080
rect 2367 990 2385 1008
rect 4311 990 4356 1026
rect 2205 576 2223 594
rect 2646 603 2673 630
rect 2718 612 2763 639
rect 3762 450 3780 468
rect 2646 189 2673 216
rect 2655 99 2754 117
rect 3069 0 3087 72
rect 4590 639 4617 666
rect 4311 450 4329 468
rect 4590 144 4617 171
rect 4311 -45 4329 -27
rect 1017 -387 1080 -306
rect 4590 -270 4617 -243
rect 4311 -486 4329 -468
rect 1008 -1035 1071 -981
rect 846 -3465 864 -3447
rect 4590 -801 4617 -774
rect 4302 -1026 4338 -990
rect 4590 -1278 4617 -1251
rect 4302 -1476 4347 -1440
rect 4590 -1773 4617 -1746
rect 4302 -1980 4347 -1935
rect 4590 -2187 4617 -2160
rect 4311 -2349 4329 -2322
rect 4590 -2718 4617 -2691
rect 4302 -2925 4347 -2889
rect 3960 -3348 4014 -3321
rect 4590 -3285 4617 -3258
rect 1035 -4599 1053 -4509
rect 4311 -3465 4329 -3447
rect 4590 -3780 4617 -3753
rect 4311 -3978 4329 -3960
rect 4590 -4194 4617 -4167
rect 4311 -4410 4329 -4392
rect 4590 -4725 4617 -4698
rect 4302 -4941 4338 -4905
rect 4590 -5220 4617 -5193
rect 4302 -5409 4347 -5382
rect 4590 -5715 4617 -5688
rect 4293 -5913 4356 -5868
rect 4590 -6129 4617 -6102
rect 4293 -6336 4338 -6300
rect 4590 -6660 4617 -6633
rect 3519 -6858 3591 -6804
<< metal1 >>
rect 4581 4806 4815 4824
rect 4581 4779 4608 4806
rect 3780 4761 4608 4779
rect 3780 4014 3798 4761
rect 4131 4707 4149 4761
rect 4284 4707 4302 4761
rect 4581 4752 4608 4761
rect 4185 4626 4203 4680
rect 4347 4626 4365 4689
rect 4653 4671 4680 4716
rect 4509 4635 4599 4662
rect 4653 4644 4707 4671
rect 4509 4626 4527 4635
rect 4185 4608 4527 4626
rect 4653 4626 4680 4644
rect 4347 4572 4365 4608
rect 4581 4563 4608 4590
rect 4131 4527 4149 4545
rect 4581 4545 4680 4563
rect 4581 4527 4617 4545
rect 4023 4509 4617 4527
rect 4023 4032 4041 4509
rect 4293 4356 4320 4374
rect 4797 4329 4815 4806
rect 4581 4311 4815 4329
rect 4581 4284 4608 4311
rect 4131 4266 4608 4284
rect 4131 4212 4149 4266
rect 4284 4212 4302 4266
rect 4581 4257 4608 4266
rect 4185 4131 4203 4185
rect 4347 4131 4365 4194
rect 4653 4176 4680 4221
rect 4509 4140 4599 4167
rect 4653 4149 4707 4176
rect 4509 4131 4527 4140
rect 4185 4113 4527 4131
rect 4653 4131 4680 4149
rect 4347 4077 4365 4113
rect 4581 4068 4608 4095
rect 4131 4032 4149 4050
rect 4581 4050 4680 4068
rect 4581 4032 4617 4050
rect 4023 4014 4617 4032
rect 2799 3996 3825 4014
rect 2799 1818 2826 3996
rect 3555 3960 3573 3996
rect 3780 3960 3798 3996
rect 3708 3879 3726 3933
rect 3618 3861 3807 3879
rect 3618 3834 3636 3861
rect 3708 3834 3726 3861
rect 3834 3834 3852 3933
rect 3564 3789 3582 3816
rect 3654 3789 3672 3816
rect 3780 3789 3798 3816
rect 4023 3789 4041 4014
rect 4797 3915 4815 4311
rect 4581 3897 4815 3915
rect 4581 3870 4608 3897
rect 3546 3771 4041 3789
rect 4131 3852 4608 3870
rect 4131 3798 4149 3852
rect 4284 3798 4302 3852
rect 4581 3843 4608 3852
rect 1836 1800 2826 1818
rect 1836 1035 1854 1800
rect 2799 1701 2826 1800
rect 4023 3618 4041 3771
rect 4185 3717 4203 3771
rect 4347 3717 4365 3780
rect 4653 3762 4680 3807
rect 4509 3726 4599 3753
rect 4653 3735 4707 3762
rect 4509 3717 4527 3726
rect 4185 3699 4527 3717
rect 4653 3717 4680 3735
rect 4347 3663 4365 3699
rect 4581 3654 4608 3681
rect 4131 3618 4149 3636
rect 4581 3636 4680 3654
rect 4581 3618 4617 3636
rect 4023 3600 4617 3618
rect 4023 3087 4041 3600
rect 4293 3528 4320 3546
rect 4797 3384 4815 3897
rect 4581 3366 4815 3384
rect 4581 3339 4608 3366
rect 4131 3321 4608 3339
rect 4131 3267 4149 3321
rect 4284 3267 4302 3321
rect 4581 3312 4608 3321
rect 4185 3186 4203 3240
rect 4347 3186 4365 3249
rect 4653 3231 4680 3276
rect 4509 3195 4599 3222
rect 4653 3204 4707 3231
rect 4509 3186 4527 3195
rect 4185 3168 4527 3186
rect 4653 3186 4680 3204
rect 4347 3132 4365 3168
rect 4581 3123 4608 3150
rect 4131 3087 4149 3105
rect 4581 3105 4680 3123
rect 4581 3087 4617 3105
rect 4023 3069 4617 3087
rect 4023 2520 4041 3069
rect 4275 2988 4320 3006
rect 4797 2817 4815 3366
rect 4581 2799 4815 2817
rect 4581 2772 4608 2799
rect 4086 2754 4608 2772
rect 4131 2700 4149 2754
rect 4284 2700 4302 2754
rect 4581 2745 4608 2754
rect 4185 2619 4203 2673
rect 4347 2619 4365 2682
rect 4653 2664 4680 2709
rect 4509 2628 4599 2655
rect 4653 2637 4707 2664
rect 4509 2619 4527 2628
rect 4185 2601 4527 2619
rect 4653 2619 4680 2637
rect 4347 2565 4365 2601
rect 4581 2556 4608 2583
rect 4131 2520 4149 2538
rect 4581 2538 4680 2556
rect 4581 2520 4617 2538
rect 4023 2502 4617 2520
rect 4023 2025 4041 2502
rect 4275 2421 4311 2439
rect 4797 2322 4815 2799
rect 4581 2304 4815 2322
rect 4581 2277 4608 2304
rect 4131 2259 4608 2277
rect 4131 2205 4149 2259
rect 4284 2205 4302 2259
rect 4581 2250 4608 2259
rect 4185 2124 4203 2178
rect 4347 2124 4365 2187
rect 4653 2169 4680 2214
rect 4509 2133 4599 2160
rect 4653 2142 4707 2169
rect 4509 2124 4527 2133
rect 4185 2106 4527 2124
rect 4653 2124 4680 2142
rect 4347 2070 4365 2106
rect 4581 2061 4608 2088
rect 4131 2025 4149 2043
rect 4581 2043 4680 2061
rect 4581 2025 4617 2043
rect 4023 2007 4617 2025
rect 4023 1782 4041 2007
rect 4275 1944 4311 1962
rect 4797 1908 4815 2304
rect 4581 1890 4815 1908
rect 4581 1863 4608 1890
rect 3978 1764 4041 1782
rect 4131 1845 4608 1863
rect 4131 1791 4149 1845
rect 4284 1791 4302 1845
rect 4581 1836 4608 1845
rect 2628 1683 2826 1701
rect 2628 1656 2655 1683
rect 2178 1638 2655 1656
rect 2178 1584 2196 1638
rect 2331 1584 2349 1638
rect 2628 1629 2655 1638
rect 2232 1503 2250 1557
rect 2394 1503 2412 1566
rect 2556 1512 2646 1539
rect 2556 1503 2574 1512
rect 2178 1476 2196 1494
rect 2232 1485 2574 1503
rect 2700 1503 2727 1593
rect 2331 1458 2349 1476
rect 2394 1449 2412 1485
rect 2628 1440 2655 1467
rect 2178 1404 2196 1422
rect 2628 1422 2727 1440
rect 2628 1404 2664 1422
rect 2088 1386 2664 1404
rect 1827 1017 1935 1035
rect 1836 972 1863 1017
rect 1908 891 1935 936
rect 2088 936 2106 1386
rect 2799 1233 2826 1683
rect 4023 1611 4041 1764
rect 4185 1710 4203 1764
rect 4347 1710 4365 1773
rect 4653 1755 4680 1800
rect 4509 1719 4599 1746
rect 4653 1728 4707 1755
rect 4509 1710 4527 1719
rect 4185 1692 4527 1710
rect 4653 1710 4680 1728
rect 4347 1656 4365 1692
rect 4581 1647 4608 1674
rect 4131 1611 4149 1629
rect 4581 1629 4680 1647
rect 4581 1611 4617 1629
rect 4023 1593 4617 1611
rect 3537 1503 3555 1521
rect 3591 1503 3618 1521
rect 2628 1215 2826 1233
rect 2628 1188 2655 1215
rect 2178 1170 2655 1188
rect 2178 1116 2196 1170
rect 2331 1116 2349 1170
rect 2628 1161 2655 1170
rect 2232 1035 2250 1089
rect 2394 1035 2412 1098
rect 2700 1080 2727 1125
rect 2556 1044 2646 1071
rect 2700 1053 2718 1080
rect 2556 1035 2574 1044
rect 2232 1017 2574 1035
rect 2700 1035 2727 1053
rect 2340 990 2367 1008
rect 2394 981 2412 1017
rect 2628 972 2655 999
rect 2178 936 2196 954
rect 2628 954 2727 972
rect 2628 936 2664 954
rect 2088 918 2664 936
rect 1908 864 1989 891
rect 1908 846 1935 864
rect 1836 783 1863 810
rect 2088 783 2106 918
rect 2799 792 2826 1215
rect 4023 1080 4041 1593
rect 4284 1503 4302 1521
rect 4347 1503 4365 1521
rect 4797 1377 4815 1890
rect 4581 1359 4815 1377
rect 4581 1332 4608 1359
rect 4131 1314 4608 1332
rect 4131 1260 4149 1314
rect 4284 1260 4302 1314
rect 4581 1305 4608 1314
rect 4185 1179 4203 1233
rect 4347 1179 4365 1242
rect 4653 1224 4680 1269
rect 4509 1188 4599 1215
rect 4653 1197 4707 1224
rect 4509 1179 4527 1188
rect 4185 1161 4527 1179
rect 4653 1179 4680 1197
rect 4347 1125 4365 1161
rect 4581 1116 4608 1143
rect 4131 1080 4149 1098
rect 4581 1098 4680 1116
rect 4581 1080 4617 1098
rect 4023 1062 4617 1080
rect 3474 1017 3510 1035
rect 3474 990 3510 999
rect 3474 936 3483 990
rect 3501 936 3510 990
rect 1710 765 2106 783
rect 2628 774 2826 792
rect 1710 459 1728 765
rect 2628 747 2655 774
rect 2070 729 2655 747
rect 2070 720 2088 729
rect 1836 702 2088 720
rect 1836 693 1872 702
rect 1845 648 1872 693
rect 2178 675 2196 729
rect 2331 675 2349 729
rect 2628 720 2655 729
rect 1917 567 1944 612
rect 2232 594 2250 648
rect 2394 594 2412 657
rect 2700 639 2727 684
rect 2556 603 2646 630
rect 2700 612 2718 639
rect 2556 594 2574 603
rect 2169 576 2205 594
rect 2232 576 2574 594
rect 2700 594 2727 612
rect 1917 540 1980 567
rect 2394 540 2412 576
rect 1917 522 1944 540
rect 2628 531 2655 558
rect 2178 495 2196 513
rect 2628 513 2727 531
rect 2628 495 2664 513
rect 1845 459 1872 486
rect 2178 477 2664 495
rect 2178 459 2196 477
rect 1710 441 2196 459
rect 1845 81 1863 441
rect 2799 378 2826 774
rect 4023 531 4041 1062
rect 4293 999 4311 1017
rect 4797 828 4815 1359
rect 4572 810 4815 828
rect 4572 783 4599 810
rect 4122 765 4599 783
rect 4122 711 4140 765
rect 4275 711 4293 765
rect 4572 756 4599 765
rect 4176 630 4194 684
rect 4338 630 4356 693
rect 4644 675 4671 720
rect 4500 639 4590 666
rect 4644 648 4698 675
rect 4500 630 4518 639
rect 4176 612 4518 630
rect 4644 630 4671 648
rect 4338 576 4356 612
rect 4572 567 4599 594
rect 4122 531 4140 549
rect 4572 549 4671 567
rect 4572 531 4608 549
rect 4014 513 4608 531
rect 3780 450 3852 468
rect 2628 360 2826 378
rect 2628 333 2655 360
rect 2178 315 2655 333
rect 2178 261 2196 315
rect 2331 261 2349 315
rect 2628 306 2655 315
rect 2232 180 2250 234
rect 2394 180 2412 243
rect 2700 225 2727 270
rect 2556 189 2646 216
rect 2700 198 2925 225
rect 2556 180 2574 189
rect 2232 162 2574 180
rect 2700 180 2727 198
rect 2394 126 2412 162
rect 2178 81 2196 99
rect 2628 99 2655 144
rect 2628 81 2664 99
rect 1845 63 2664 81
rect 1035 -306 1053 -63
rect 936 -486 945 -468
rect 963 -486 1062 -468
rect 1071 -1017 1188 -990
rect 1188 -1449 1251 -1440
rect 1188 -1467 1206 -1449
rect 1188 -1476 1251 -1467
rect 2907 -3321 2925 198
rect 4014 45 4032 513
rect 4284 450 4311 468
rect 4797 333 4815 810
rect 4572 315 4815 333
rect 4572 288 4599 315
rect 4122 270 4599 288
rect 4122 216 4140 270
rect 4275 216 4293 270
rect 4572 261 4599 270
rect 4176 135 4194 189
rect 4338 135 4356 198
rect 4644 180 4671 225
rect 4500 144 4590 171
rect 4644 153 4698 180
rect 4500 135 4518 144
rect 4176 117 4518 135
rect 4644 135 4671 153
rect 4338 81 4356 117
rect 3087 36 4032 45
rect 4572 72 4599 99
rect 4122 36 4140 54
rect 4572 54 4671 72
rect 4572 36 4608 54
rect 3087 18 4608 36
rect 4014 -378 4032 18
rect 4293 -45 4311 -27
rect 4797 -81 4815 315
rect 4572 -99 4815 -81
rect 4572 -126 4599 -99
rect 4122 -144 4599 -126
rect 4122 -198 4140 -144
rect 4275 -198 4293 -144
rect 4572 -153 4599 -144
rect 4176 -279 4194 -225
rect 4338 -279 4356 -216
rect 4644 -234 4671 -189
rect 4500 -270 4590 -243
rect 4644 -261 4698 -234
rect 4500 -279 4518 -270
rect 4176 -297 4518 -279
rect 4644 -279 4671 -261
rect 4338 -333 4356 -297
rect 4572 -342 4599 -315
rect 4122 -378 4140 -360
rect 4572 -360 4671 -342
rect 4572 -378 4608 -360
rect 4014 -396 4608 -378
rect 4014 -909 4032 -396
rect 4275 -486 4311 -468
rect 4797 -612 4815 -99
rect 4572 -630 4815 -612
rect 4572 -657 4599 -630
rect 4122 -675 4599 -657
rect 4122 -729 4140 -675
rect 4275 -729 4293 -675
rect 4572 -684 4599 -675
rect 4176 -810 4194 -756
rect 4338 -810 4356 -747
rect 4644 -765 4671 -720
rect 4500 -801 4590 -774
rect 4644 -792 4698 -765
rect 4500 -810 4518 -801
rect 4176 -828 4518 -810
rect 4644 -810 4671 -792
rect 4338 -864 4356 -828
rect 4572 -873 4599 -846
rect 4122 -909 4140 -891
rect 4572 -891 4671 -873
rect 4572 -909 4608 -891
rect 4014 -927 4608 -909
rect 4014 -1386 4032 -927
rect 4275 -1017 4302 -999
rect 4797 -1089 4815 -630
rect 4572 -1107 4815 -1089
rect 4572 -1134 4599 -1107
rect 4122 -1152 4599 -1134
rect 4122 -1206 4140 -1152
rect 4275 -1206 4293 -1152
rect 4572 -1161 4599 -1152
rect 4176 -1287 4194 -1233
rect 4338 -1287 4356 -1224
rect 4644 -1242 4671 -1197
rect 4500 -1278 4590 -1251
rect 4644 -1269 4698 -1242
rect 4500 -1287 4518 -1278
rect 4176 -1305 4518 -1287
rect 4644 -1287 4671 -1269
rect 4338 -1341 4356 -1305
rect 4572 -1350 4599 -1323
rect 4122 -1386 4140 -1368
rect 4572 -1368 4671 -1350
rect 4572 -1386 4608 -1368
rect 4014 -1404 4608 -1386
rect 3717 -1935 3735 -1863
rect 4014 -1881 4032 -1404
rect 4293 -1467 4302 -1449
rect 4797 -1584 4815 -1107
rect 4572 -1602 4815 -1584
rect 4572 -1629 4599 -1602
rect 4122 -1647 4599 -1629
rect 4122 -1701 4140 -1647
rect 4275 -1701 4293 -1647
rect 4572 -1656 4599 -1647
rect 4176 -1782 4194 -1728
rect 4338 -1782 4356 -1719
rect 4644 -1737 4671 -1692
rect 4500 -1773 4590 -1746
rect 4644 -1764 4698 -1737
rect 4500 -1782 4518 -1773
rect 4176 -1800 4518 -1782
rect 4644 -1782 4671 -1764
rect 4338 -1836 4356 -1800
rect 4572 -1845 4599 -1818
rect 4122 -1881 4140 -1863
rect 4572 -1863 4671 -1845
rect 4572 -1881 4608 -1863
rect 4014 -1899 4608 -1881
rect 4014 -2295 4032 -1899
rect 4266 -1962 4302 -1944
rect 4347 -1962 4356 -1944
rect 4797 -1998 4815 -1602
rect 4572 -2016 4815 -1998
rect 4572 -2043 4599 -2016
rect 4122 -2061 4599 -2043
rect 4122 -2115 4140 -2061
rect 4275 -2115 4293 -2061
rect 4572 -2070 4599 -2061
rect 4176 -2196 4194 -2142
rect 4338 -2196 4356 -2133
rect 4644 -2151 4671 -2106
rect 4500 -2187 4590 -2160
rect 4644 -2178 4698 -2151
rect 4500 -2196 4518 -2187
rect 4176 -2214 4518 -2196
rect 4644 -2196 4671 -2178
rect 4338 -2250 4356 -2214
rect 4572 -2259 4599 -2232
rect 4122 -2295 4140 -2277
rect 4572 -2277 4671 -2259
rect 4572 -2295 4608 -2277
rect 4014 -2313 4608 -2295
rect 3564 -2349 3582 -2331
rect 3600 -2367 3618 -2349
rect 3564 -2385 3582 -2367
rect 4014 -2826 4032 -2313
rect 4797 -2529 4815 -2016
rect 4572 -2547 4815 -2529
rect 4572 -2574 4599 -2547
rect 4122 -2592 4599 -2574
rect 4122 -2646 4140 -2592
rect 4275 -2646 4293 -2592
rect 4572 -2601 4599 -2592
rect 4176 -2727 4194 -2673
rect 4338 -2727 4356 -2664
rect 4644 -2682 4671 -2637
rect 4500 -2718 4590 -2691
rect 4644 -2709 4698 -2682
rect 4500 -2727 4518 -2718
rect 4176 -2745 4518 -2727
rect 4644 -2727 4671 -2709
rect 4338 -2781 4356 -2745
rect 4572 -2790 4599 -2763
rect 4122 -2826 4140 -2808
rect 4572 -2808 4671 -2790
rect 4572 -2826 4608 -2808
rect 4014 -2844 4608 -2826
rect 3465 -2916 3483 -2898
rect 3501 -2916 3510 -2898
rect 2907 -3348 3960 -3321
rect 4041 -3393 4059 -2844
rect 4257 -2916 4302 -2898
rect 4788 -3096 4806 -2547
rect 4572 -3114 4806 -3096
rect 4572 -3141 4599 -3114
rect 4122 -3159 4599 -3141
rect 4122 -3213 4140 -3159
rect 4275 -3213 4293 -3159
rect 4572 -3168 4599 -3159
rect 4176 -3294 4194 -3240
rect 4338 -3294 4356 -3231
rect 4644 -3249 4671 -3204
rect 4500 -3285 4590 -3258
rect 4644 -3276 4698 -3249
rect 4500 -3294 4518 -3285
rect 4176 -3312 4518 -3294
rect 4644 -3294 4671 -3276
rect 4338 -3348 4356 -3312
rect 4572 -3357 4599 -3330
rect 4122 -3393 4140 -3375
rect 4572 -3375 4671 -3357
rect 4572 -3393 4608 -3375
rect 4014 -3411 4608 -3393
rect 864 -3465 927 -3447
rect 4014 -3888 4032 -3411
rect 4275 -3465 4311 -3447
rect 4788 -3591 4806 -3114
rect 4572 -3609 4806 -3591
rect 4572 -3636 4599 -3609
rect 4122 -3654 4599 -3636
rect 4122 -3708 4140 -3654
rect 4275 -3708 4293 -3654
rect 4572 -3663 4599 -3654
rect 4176 -3789 4194 -3735
rect 4338 -3789 4356 -3726
rect 4644 -3744 4671 -3699
rect 4500 -3780 4590 -3753
rect 4644 -3771 4698 -3744
rect 4500 -3789 4518 -3780
rect 4176 -3807 4518 -3789
rect 4644 -3789 4671 -3771
rect 4338 -3843 4356 -3807
rect 4572 -3852 4599 -3825
rect 4122 -3888 4140 -3870
rect 4572 -3870 4671 -3852
rect 4572 -3888 4608 -3870
rect 4014 -3906 4608 -3888
rect 4014 -4302 4032 -3906
rect 4284 -3978 4311 -3960
rect 4788 -4005 4806 -3609
rect 4572 -4023 4806 -4005
rect 4572 -4050 4599 -4023
rect 4122 -4068 4599 -4050
rect 4122 -4122 4140 -4068
rect 4275 -4122 4293 -4068
rect 4572 -4077 4599 -4068
rect 4176 -4203 4194 -4149
rect 4338 -4203 4356 -4140
rect 4644 -4158 4671 -4113
rect 4500 -4194 4590 -4167
rect 4644 -4185 4698 -4158
rect 4500 -4203 4518 -4194
rect 4176 -4221 4518 -4203
rect 4644 -4203 4671 -4185
rect 4338 -4257 4356 -4221
rect 4572 -4266 4599 -4239
rect 4122 -4302 4140 -4284
rect 4572 -4284 4671 -4266
rect 4572 -4302 4608 -4284
rect 4014 -4320 4608 -4302
rect 972 -4410 1035 -4392
rect 1035 -4905 1053 -4599
rect 4014 -4833 4032 -4320
rect 4275 -4410 4311 -4392
rect 4788 -4536 4806 -4023
rect 4572 -4554 4806 -4536
rect 4572 -4581 4599 -4554
rect 4122 -4599 4599 -4581
rect 4122 -4653 4140 -4599
rect 4275 -4653 4293 -4599
rect 4572 -4608 4599 -4599
rect 4176 -4734 4194 -4680
rect 4338 -4734 4356 -4671
rect 4644 -4689 4671 -4644
rect 4500 -4725 4590 -4698
rect 4644 -4716 4698 -4689
rect 4500 -4734 4518 -4725
rect 4176 -4752 4518 -4734
rect 4644 -4734 4671 -4716
rect 4338 -4788 4356 -4752
rect 4572 -4797 4599 -4770
rect 4122 -4833 4140 -4815
rect 4572 -4815 4671 -4797
rect 4572 -4833 4608 -4815
rect 4014 -4851 4608 -4833
rect 1152 -5364 1179 -5274
rect 4014 -5328 4032 -4851
rect 4239 -4932 4302 -4914
rect 4788 -5031 4806 -4554
rect 4572 -5049 4806 -5031
rect 4572 -5076 4599 -5049
rect 4122 -5094 4599 -5076
rect 4122 -5148 4140 -5094
rect 4275 -5148 4293 -5094
rect 4572 -5103 4599 -5094
rect 4176 -5229 4194 -5175
rect 4338 -5229 4356 -5166
rect 4644 -5184 4671 -5139
rect 4500 -5220 4590 -5193
rect 4644 -5211 4698 -5184
rect 4500 -5229 4518 -5220
rect 4176 -5247 4518 -5229
rect 4644 -5229 4671 -5211
rect 4338 -5283 4356 -5247
rect 4572 -5292 4599 -5265
rect 4122 -5328 4140 -5310
rect 4572 -5310 4635 -5292
rect 4572 -5328 4608 -5310
rect 4014 -5346 4608 -5328
rect 4014 -5823 4032 -5346
rect 4275 -5400 4302 -5382
rect 4788 -5526 4806 -5049
rect 4572 -5544 4806 -5526
rect 4572 -5571 4599 -5544
rect 4122 -5589 4599 -5571
rect 4122 -5643 4140 -5589
rect 4275 -5643 4293 -5589
rect 4572 -5598 4599 -5589
rect 4176 -5724 4194 -5670
rect 4338 -5724 4356 -5661
rect 4644 -5679 4671 -5634
rect 4500 -5715 4590 -5688
rect 4644 -5706 4698 -5679
rect 4500 -5724 4518 -5715
rect 4176 -5742 4518 -5724
rect 4644 -5724 4671 -5706
rect 4338 -5778 4356 -5742
rect 4572 -5787 4599 -5760
rect 4122 -5823 4140 -5805
rect 4572 -5805 4671 -5787
rect 4572 -5823 4608 -5805
rect 4014 -5841 4608 -5823
rect 3753 -5904 3771 -5877
rect 4014 -6237 4032 -5841
rect 4257 -5895 4293 -5877
rect 4788 -5940 4806 -5544
rect 4572 -5958 4806 -5940
rect 4572 -5985 4599 -5958
rect 4122 -6003 4599 -5985
rect 4122 -6057 4140 -6003
rect 4275 -6057 4293 -6003
rect 4572 -6012 4599 -6003
rect 4176 -6138 4194 -6084
rect 4338 -6138 4356 -6075
rect 4644 -6093 4671 -6048
rect 4500 -6129 4590 -6102
rect 4644 -6120 4698 -6093
rect 4500 -6138 4518 -6129
rect 4176 -6156 4518 -6138
rect 4644 -6138 4671 -6120
rect 4338 -6192 4356 -6156
rect 4572 -6201 4599 -6174
rect 4122 -6237 4140 -6219
rect 4572 -6219 4671 -6201
rect 4572 -6237 4608 -6219
rect 4014 -6255 4608 -6237
rect 4014 -6768 4032 -6255
rect 4266 -6327 4293 -6309
rect 4788 -6471 4806 -5958
rect 4572 -6489 4806 -6471
rect 4572 -6516 4599 -6489
rect 4122 -6534 4599 -6516
rect 4122 -6588 4140 -6534
rect 4275 -6588 4293 -6534
rect 4572 -6543 4599 -6534
rect 4176 -6669 4194 -6615
rect 4338 -6669 4356 -6606
rect 4644 -6624 4671 -6579
rect 4500 -6660 4590 -6633
rect 4644 -6651 4698 -6624
rect 4500 -6669 4518 -6660
rect 4176 -6687 4518 -6669
rect 4644 -6669 4671 -6651
rect 4338 -6723 4356 -6687
rect 4572 -6732 4599 -6705
rect 4122 -6768 4140 -6750
rect 4572 -6750 4671 -6732
rect 4572 -6768 4608 -6750
rect 4014 -6786 4608 -6768
rect 3456 -6840 3474 -6822
rect 3501 -6840 3519 -6822
<< m2contact >>
rect 4248 4356 4293 4374
rect 4185 2988 4275 3006
rect 2133 1476 2178 1494
rect 3618 1494 3708 1530
rect 1989 864 2016 891
rect 4095 1503 4284 1521
rect 3438 999 3537 1017
rect 2133 576 2169 594
rect 4212 990 4293 1026
rect 3852 450 3924 468
rect 1035 -63 1053 36
rect 1062 -486 1134 -468
rect 1188 -1017 1350 -990
rect 1206 -1467 1269 -1449
rect 4239 450 4284 468
rect 4212 -45 4293 -27
rect 4212 -486 4275 -468
rect 4185 -1035 4275 -990
rect 4221 -1476 4293 -1440
rect 3699 -1980 3762 -1935
rect 4203 -1971 4266 -1935
rect 3618 -2367 3681 -2349
rect 4293 -2367 4329 -2349
rect 3510 -2916 3546 -2898
rect 4176 -2925 4257 -2889
rect 927 -3465 981 -3447
rect 4230 -3465 4275 -3447
rect 4212 -3978 4284 -3960
rect 1035 -4410 1107 -4392
rect 4131 -4410 4275 -4392
rect 999 -4950 1080 -4905
rect 1152 -5427 1179 -5364
rect 4149 -4941 4239 -4905
rect 4185 -5418 4275 -5382
rect 3771 -5913 3843 -5868
rect 4176 -5904 4257 -5868
<< metal2 >>
rect 666 4356 4248 4374
rect 666 -207 693 4356
rect 1035 2988 4185 3006
rect 1035 36 1053 2988
rect 3708 1503 4095 1521
rect 1998 1476 2133 1494
rect 1998 891 2016 1476
rect 3537 999 4212 1017
rect 2016 864 2070 891
rect 2052 594 2070 864
rect 2052 576 2133 594
rect 3924 450 4239 468
rect 3888 -45 4212 -27
rect 3888 -207 3906 -45
rect 666 -243 3906 -207
rect 666 -3960 693 -243
rect 1134 -486 4212 -468
rect 3654 -990 3744 -981
rect 1350 -999 3744 -990
rect 1350 -1017 4185 -999
rect 3654 -1035 3744 -1017
rect 1269 -1467 4221 -1449
rect 3690 -1962 3699 -1944
rect 3762 -1962 4203 -1944
rect 3681 -2367 4293 -2349
rect 3546 -2916 4176 -2898
rect 981 -3465 4230 -3447
rect 666 -3978 4212 -3960
rect 1107 -4410 4131 -4392
rect 1080 -4932 4149 -4914
rect 1125 -5400 1152 -5382
rect 1179 -5400 4185 -5382
rect 3843 -5895 4176 -5877
<< m123contact >>
rect 4221 3528 4293 3546
rect 4158 2412 4275 2448
rect 4203 1935 4275 1962
rect 3555 1494 3591 1539
rect 2295 1458 2331 1476
rect 2286 990 2340 1008
rect 3483 918 3501 990
rect 1980 540 2034 567
rect 945 -486 963 -468
rect 1134 -1494 1188 -1431
rect 3708 -1863 3753 -1800
rect 3564 -2367 3600 -2349
rect 3483 -2934 3501 -2889
rect 936 -4419 972 -4383
rect 1134 -5274 1197 -5211
rect 3690 -5913 3753 -5868
rect 4203 -6327 4266 -6309
rect 3474 -6858 3501 -6813
<< metal3 >>
rect 945 3528 4221 3546
rect 945 -468 963 3528
rect 945 -4383 963 -486
rect 1152 2421 4158 2439
rect 1152 -1431 1179 2421
rect 3717 1944 4203 1962
rect 2295 1296 2313 1458
rect 2016 1278 2313 1296
rect 2016 909 2034 1278
rect 2286 909 2304 990
rect 2016 891 2304 909
rect 2016 567 2034 891
rect 1152 -5211 1179 -1494
rect 3483 -2889 3501 918
rect 3483 -6813 3501 -2934
rect 3564 -2349 3582 1494
rect 3717 -1800 3735 1944
rect 3564 -6309 3582 -2367
rect 3717 -5868 3735 -1863
rect 3564 -6327 4203 -6309
<< labels >>
rlabel polysilicon 1746 945 1746 945 1 s0
rlabel polysilicon 1800 549 1800 549 1 s1
rlabel metal1 1845 1341 1845 1341 1 vdd
rlabel metal1 1962 72 1962 72 1 gnd
rlabel metal1 2745 207 2745 207 1 D3
rlabel polycontact 2745 621 2745 621 1 D2
rlabel polycontact 2727 1062 2727 1062 1 D1
rlabel polycontact 2736 1539 2736 1539 1 D0
rlabel metal1 1962 873 1962 873 1 s0_not
rlabel metal1 1971 549 1971 549 1 s1_not
rlabel metal1 4671 -4707 4671 -4707 1 and_a0
rlabel metal1 4671 -4176 4671 -4176 1 and_a1
rlabel metal1 4671 -3762 4671 -3762 1 and_a2
rlabel metal1 4680 -3258 4680 -3258 1 and_a3
rlabel metal1 4671 -6642 4671 -6642 1 and_b0
rlabel metal1 4680 -6111 4680 -6111 1 and_b1
rlabel metal1 4689 -5697 4689 -5697 1 and_b2
rlabel metal1 4680 -5202 4680 -5202 1 and_b3
rlabel metal1 4680 657 4680 657 1 comp_a3
rlabel metal1 4680 171 4680 171 1 comp_a2
rlabel metal1 4680 -243 4680 -243 1 comp_a1
rlabel metal1 4680 -783 4680 -783 1 comp_a0
rlabel metal1 4671 -1260 4671 -1260 1 comp_b3
rlabel metal1 4680 -1755 4680 -1755 1 comp_b2
rlabel metal1 4680 -2160 4680 -2160 1 comp_b1
rlabel metal1 4680 -2700 4680 -2700 1 comp_b0
rlabel metal1 4689 1215 4689 1215 1 adsub_b0
rlabel metal1 4680 1746 4680 1746 1 adsub_b1
rlabel polysilicon 4329 1674 4329 1674 1 b1
rlabel metal1 4689 2160 4689 2160 1 adsub_b2
rlabel polysilicon 4329 2088 4329 2088 1 b2
rlabel metal1 4689 2646 4689 2646 1 adsub_b3
rlabel polysilicon 4329 2592 4329 2592 1 b3
rlabel polysilicon 4329 3150 4329 3150 1 a0
rlabel metal1 4689 3213 4689 3213 1 adsub_a0
rlabel metal1 4689 3744 4689 3744 1 adsub_a1
rlabel metal1 4689 4158 4689 4158 1 adsub_a2
rlabel metal1 4680 4662 4680 4662 1 adsub_a3
rlabel polysilicon 4329 4599 4329 4599 1 a3
rlabel polysilicon 4329 4095 4329 4095 1 a2
rlabel polysilicon 4329 3681 4329 3681 1 a1
rlabel polysilicon 3942 3870 3942 3870 1 D
rlabel polysilicon 4329 1143 4329 1143 1 b0
<< end >>
