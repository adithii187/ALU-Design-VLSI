magic
tech scmos
magscale 9 1
timestamp 1698857296
<< nwell >>
rect -19 1 56 13
<< ntransistor >>
rect -12 -24 -10 -18
rect 7 -24 9 -18
rect 29 -24 31 -18
rect 47 -24 49 -18
<< ptransistor >>
rect -12 4 -10 11
rect 7 4 9 11
rect 29 4 31 11
rect 47 4 49 11
<< ndiffusion >>
rect -18 -19 -12 -18
rect -18 -23 -17 -19
rect -13 -23 -12 -19
rect -18 -24 -12 -23
rect -10 -19 -4 -18
rect -10 -23 -9 -19
rect -5 -23 -4 -19
rect -10 -24 -4 -23
rect 1 -19 7 -18
rect 1 -23 2 -19
rect 6 -23 7 -19
rect 1 -24 7 -23
rect 9 -19 15 -18
rect 9 -23 10 -19
rect 14 -23 15 -19
rect 9 -24 15 -23
rect 22 -19 29 -18
rect 22 -23 23 -19
rect 27 -23 29 -19
rect 22 -24 29 -23
rect 31 -19 37 -18
rect 31 -23 32 -19
rect 36 -23 37 -19
rect 31 -24 37 -23
rect 40 -19 47 -18
rect 40 -23 41 -19
rect 45 -23 47 -19
rect 40 -24 47 -23
rect 49 -19 55 -18
rect 49 -23 50 -19
rect 54 -23 55 -19
rect 49 -24 55 -23
<< pdiffusion >>
rect -18 9 -12 11
rect -18 5 -17 9
rect -13 5 -12 9
rect -18 4 -12 5
rect -10 9 -4 11
rect -10 5 -9 9
rect -5 5 -4 9
rect -10 4 -4 5
rect 1 9 7 11
rect 1 5 2 9
rect 6 5 7 9
rect 1 4 7 5
rect 9 9 15 11
rect 9 5 10 9
rect 14 5 15 9
rect 9 4 15 5
rect 22 9 29 11
rect 22 5 23 9
rect 27 5 29 9
rect 22 4 29 5
rect 31 9 37 11
rect 31 5 32 9
rect 36 5 37 9
rect 31 4 37 5
rect 40 9 47 11
rect 40 5 41 9
rect 45 5 47 9
rect 40 4 47 5
rect 49 9 55 11
rect 49 5 50 9
rect 54 5 55 9
rect 49 4 55 5
<< ndcontact >>
rect -17 -23 -13 -19
rect -9 -23 -5 -19
rect 2 -23 6 -19
rect 10 -23 14 -19
rect 23 -23 27 -19
rect 32 -23 36 -19
rect 41 -23 45 -19
rect 50 -23 54 -19
<< pdcontact >>
rect -17 5 -13 9
rect -9 5 -5 9
rect 2 5 6 9
rect 10 5 14 9
rect 23 5 27 9
rect 32 5 36 9
rect 41 5 45 9
rect 50 5 54 9
<< psubstratepcontact >>
rect 27 -37 31 -33
rect 37 -37 41 -33
<< nsubstratencontact >>
rect 27 18 31 22
rect 37 18 41 22
<< polysilicon >>
rect -24 17 9 19
rect -24 -28 -22 17
rect -12 11 -10 14
rect 7 11 9 17
rect 29 11 31 16
rect 47 11 49 16
rect -12 -13 -10 4
rect 7 0 9 4
rect 29 -6 31 4
rect 47 -6 49 4
rect 26 -10 31 -6
rect 42 -10 49 -6
rect -12 -15 9 -13
rect -12 -18 -10 -17
rect 7 -18 9 -15
rect 29 -18 31 -10
rect 47 -18 49 -10
rect -12 -28 -10 -24
rect -24 -30 -10 -28
rect -12 -45 -10 -30
rect 7 -40 9 -24
rect 29 -31 31 -24
rect 47 -40 49 -24
rect 7 -42 49 -40
rect 61 -45 63 -6
rect -12 -47 63 -45
<< polycontact >>
rect 22 -10 26 -6
rect 57 -10 61 -6
<< metal1 >>
rect -17 25 21 29
rect -17 9 -13 25
rect -17 -19 -13 5
rect -9 20 14 24
rect -9 9 -5 20
rect 10 9 14 20
rect -9 -19 -5 5
rect 2 -19 6 5
rect 10 -19 14 5
rect 17 -6 21 25
rect 23 9 27 22
rect 31 18 37 22
rect 41 9 45 22
rect 17 -10 22 -6
rect 32 -12 36 5
rect 17 -16 36 -12
rect 2 -33 6 -23
rect 17 -33 21 -16
rect 32 -19 36 -16
rect 50 -6 54 5
rect 50 -10 57 -6
rect 50 -19 54 -10
rect 2 -37 21 -33
rect 23 -37 27 -23
rect 31 -37 37 -33
rect 41 -37 45 -23
<< labels >>
rlabel polysilicon 27 -9 27 -9 1 va
rlabel metal1 35 -8 35 -8 1 vab
rlabel polysilicon 45 -8 45 -8 1 vb
rlabel metal1 53 -8 53 -8 1 vbb
rlabel metal1 34 19 34 19 5 vdd
rlabel metal1 34 -35 34 -35 1 gnd
rlabel metal1 3 22 3 22 1 vout
<< end >>
