magic
tech scmos
timestamp 1700736304
<< nwell >>
rect 4662 6201 4851 6255
rect 4194 6048 4518 6138
rect 4662 6093 4815 6201
rect 4662 6084 4725 6093
rect 4743 6084 4815 6093
rect 4662 5706 4851 5760
rect 4194 5553 4518 5643
rect 4662 5598 4815 5706
rect 4662 5589 4725 5598
rect 4743 5589 4815 5598
rect 4662 5292 4851 5346
rect 4194 5139 4518 5229
rect 4662 5184 4815 5292
rect 4662 5175 4725 5184
rect 4743 5175 4815 5184
rect 4662 4761 4851 4815
rect 4194 4608 4518 4698
rect 4662 4653 4815 4761
rect 4662 4644 4725 4653
rect 4743 4644 4815 4653
rect 4662 3762 4851 3816
rect 4194 3609 4518 3699
rect 4662 3654 4815 3762
rect 4662 3645 4725 3654
rect 4743 3645 4815 3654
rect 4662 3267 4851 3321
rect 4194 3114 4518 3204
rect 4662 3159 4815 3267
rect 4662 3150 4725 3159
rect 4743 3150 4815 3159
rect 3636 2871 3987 2988
rect 4662 2853 4851 2907
rect 4194 2700 4518 2790
rect 4662 2745 4815 2853
rect 4662 2736 4725 2745
rect 4743 2736 4815 2745
rect 4662 2322 4851 2376
rect 4194 2169 4518 2259
rect 4662 2214 4815 2322
rect 4662 2205 4725 2214
rect 4743 2205 4815 2214
rect 2988 1710 3168 1764
rect 5463 1719 5652 1773
rect 2520 1557 2844 1647
rect 2988 1602 3141 1710
rect 2988 1593 3051 1602
rect 3069 1593 3141 1602
rect 4995 1566 5319 1656
rect 5463 1611 5616 1719
rect 5463 1602 5526 1611
rect 5544 1602 5616 1611
rect 2988 1242 3168 1296
rect 2187 1071 2376 1098
rect 2520 1089 2844 1179
rect 2988 1134 3141 1242
rect 5463 1224 5652 1278
rect 2988 1125 3051 1134
rect 3069 1125 3141 1134
rect 4995 1071 5319 1161
rect 5463 1116 5616 1224
rect 5463 1107 5526 1116
rect 5544 1107 5616 1116
rect 2187 1053 2214 1071
rect 2322 1053 2376 1071
rect 2196 945 2349 1053
rect 2196 936 2259 945
rect 2277 936 2349 945
rect 2988 801 3168 855
rect 5463 810 5652 864
rect 2196 729 2385 774
rect 2205 621 2358 729
rect 2520 648 2844 738
rect 2988 693 3141 801
rect 2988 684 3051 693
rect 3069 684 3141 693
rect 4995 657 5319 747
rect 5463 702 5616 810
rect 5463 693 5526 702
rect 5544 693 5616 702
rect 2205 612 2268 621
rect 2286 612 2358 621
rect 2988 387 3177 441
rect 2520 234 2844 324
rect 2988 279 3141 387
rect 2988 270 3051 279
rect 3069 270 3141 279
rect 5463 279 5652 333
rect 4995 126 5319 216
rect 5463 171 5616 279
rect 5463 162 5526 171
rect 5544 162 5616 171
rect 3852 -90 4041 -36
rect 6642 -45 6831 9
rect 3384 -243 3708 -153
rect 3852 -198 4005 -90
rect 6174 -198 6498 -108
rect 6642 -153 6795 -45
rect 6642 -162 6705 -153
rect 6723 -162 6795 -153
rect 3852 -207 3915 -198
rect 3933 -207 4005 -198
rect 3852 -585 4041 -531
rect 6642 -540 6831 -486
rect 3384 -738 3708 -648
rect 3852 -693 4005 -585
rect 6174 -693 6498 -603
rect 6642 -648 6795 -540
rect 6642 -657 6705 -648
rect 6723 -657 6795 -648
rect 3852 -702 3915 -693
rect 3933 -702 4005 -693
rect 3852 -999 4041 -945
rect 6642 -954 6831 -900
rect 3384 -1152 3708 -1062
rect 3852 -1107 4005 -999
rect 6174 -1107 6498 -1017
rect 6642 -1062 6795 -954
rect 6642 -1071 6705 -1062
rect 6723 -1071 6795 -1062
rect 3852 -1116 3915 -1107
rect 3933 -1116 4005 -1107
rect 3852 -1530 4041 -1476
rect 6642 -1485 6831 -1431
rect 3384 -1683 3708 -1593
rect 3852 -1638 4005 -1530
rect 6174 -1638 6498 -1548
rect 6642 -1593 6795 -1485
rect 6642 -1602 6705 -1593
rect 6723 -1602 6795 -1593
rect 3852 -1647 3915 -1638
rect 3933 -1647 4005 -1638
rect 5517 -2241 5706 -2187
rect 3807 -2358 3996 -2304
rect 3339 -2511 3663 -2421
rect 3807 -2466 3960 -2358
rect 5049 -2394 5373 -2304
rect 5517 -2349 5670 -2241
rect 5517 -2358 5580 -2349
rect 5598 -2358 5670 -2349
rect 3807 -2475 3870 -2466
rect 3888 -2475 3960 -2466
rect 5517 -2718 5706 -2664
rect 3807 -2853 3996 -2799
rect 3339 -3006 3663 -2916
rect 3807 -2961 3960 -2853
rect 5049 -2871 5373 -2781
rect 5517 -2826 5670 -2718
rect 5517 -2835 5580 -2826
rect 5598 -2835 5670 -2826
rect 3807 -2970 3870 -2961
rect 3888 -2970 3960 -2961
rect 5517 -3114 5706 -3060
rect 3807 -3267 3996 -3213
rect 5049 -3267 5373 -3177
rect 5517 -3222 5670 -3114
rect 5517 -3231 5580 -3222
rect 5598 -3231 5670 -3222
rect 3339 -3420 3663 -3330
rect 3807 -3375 3960 -3267
rect 3807 -3384 3870 -3375
rect 3888 -3384 3960 -3375
rect 5517 -3582 5706 -3528
rect 5049 -3735 5373 -3645
rect 5517 -3690 5670 -3582
rect 5517 -3699 5580 -3690
rect 5598 -3699 5670 -3690
rect 3807 -3798 3996 -3744
rect 3339 -3951 3663 -3861
rect 3807 -3906 3960 -3798
rect 3807 -3915 3870 -3906
rect 3888 -3915 3960 -3906
<< ntransistor >>
rect 4725 6003 4743 6030
rect 4266 5949 4284 5976
rect 4428 5949 4446 5976
rect 4725 5508 4743 5535
rect 4266 5454 4284 5481
rect 4428 5454 4446 5481
rect 4725 5094 4743 5121
rect 4266 5040 4284 5067
rect 4428 5040 4446 5067
rect 4725 4563 4743 4590
rect 4266 4509 4284 4536
rect 4428 4509 4446 4536
rect 4725 3564 4743 3591
rect 4266 3510 4284 3537
rect 4428 3510 4446 3537
rect 4725 3069 4743 3096
rect 4266 3015 4284 3042
rect 4428 3015 4446 3042
rect 3699 2772 3717 2799
rect 3789 2772 3807 2799
rect 3915 2772 3933 2799
rect 3051 1512 3069 1539
rect 2592 1458 2610 1485
rect 2754 1458 2772 1485
rect 4725 2655 4743 2682
rect 4266 2601 4284 2628
rect 4428 2601 4446 2628
rect 4725 2124 4743 2151
rect 4266 2070 4284 2097
rect 4428 2070 4446 2097
rect 3051 1044 3069 1071
rect 5526 1521 5544 1548
rect 5067 1467 5085 1494
rect 5229 1467 5247 1494
rect 2592 990 2610 1017
rect 2754 990 2772 1017
rect 2259 855 2277 882
rect 5526 1026 5544 1053
rect 5067 972 5085 999
rect 5229 972 5247 999
rect 3051 603 3069 630
rect 2268 531 2286 558
rect 2592 549 2610 576
rect 2727 549 2745 576
rect 2754 549 2772 576
rect 3051 189 3069 216
rect 2592 135 2610 162
rect 2709 135 2727 162
rect 2754 135 2772 162
rect 3915 -288 3933 -261
rect 3456 -342 3474 -315
rect 3618 -342 3636 -315
rect 3915 -783 3933 -756
rect 3456 -837 3474 -810
rect 3618 -837 3636 -810
rect 3915 -1197 3933 -1170
rect 3456 -1251 3474 -1224
rect 3618 -1251 3636 -1224
rect 3915 -1728 3933 -1701
rect 3456 -1782 3474 -1755
rect 3618 -1782 3636 -1755
rect 3870 -2556 3888 -2529
rect 3411 -2610 3429 -2583
rect 3573 -2610 3591 -2583
rect 5526 612 5544 639
rect 5067 558 5085 585
rect 5229 558 5247 585
rect 5526 81 5544 108
rect 5067 27 5085 54
rect 5229 27 5247 54
rect 6705 -243 6723 -216
rect 6246 -297 6264 -270
rect 6408 -297 6426 -270
rect 6705 -738 6723 -711
rect 6246 -792 6264 -765
rect 6408 -792 6426 -765
rect 6705 -1152 6723 -1125
rect 6246 -1206 6264 -1179
rect 6408 -1206 6426 -1179
rect 6705 -1683 6723 -1656
rect 6246 -1737 6264 -1710
rect 6408 -1737 6426 -1710
rect 5580 -2439 5598 -2412
rect 5121 -2493 5139 -2466
rect 5283 -2493 5301 -2466
rect 5580 -2916 5598 -2889
rect 5121 -2970 5139 -2943
rect 5283 -2970 5301 -2943
rect 3870 -3051 3888 -3024
rect 3411 -3105 3429 -3078
rect 3573 -3105 3591 -3078
rect 5580 -3312 5598 -3285
rect 5121 -3366 5139 -3339
rect 5283 -3366 5301 -3339
rect 3870 -3465 3888 -3438
rect 3411 -3519 3429 -3492
rect 3573 -3519 3591 -3492
rect 5580 -3780 5598 -3753
rect 5121 -3834 5139 -3807
rect 5283 -3834 5301 -3807
rect 3870 -3996 3888 -3969
rect 3411 -4050 3429 -4023
rect 3573 -4050 3591 -4023
<< ptransistor >>
rect 4266 6075 4284 6120
rect 4428 6075 4446 6120
rect 4725 6102 4743 6156
rect 4266 5580 4284 5625
rect 4428 5580 4446 5625
rect 4725 5607 4743 5661
rect 4266 5166 4284 5211
rect 4428 5166 4446 5211
rect 4725 5193 4743 5247
rect 4266 4635 4284 4680
rect 4428 4635 4446 4680
rect 4725 4662 4743 4716
rect 4266 3636 4284 3681
rect 4428 3636 4446 3681
rect 4725 3663 4743 3717
rect 4266 3141 4284 3186
rect 4428 3141 4446 3186
rect 4725 3168 4743 3222
rect 3699 2889 3717 2934
rect 3789 2889 3807 2934
rect 3915 2889 3933 2934
rect 2592 1584 2610 1629
rect 2754 1584 2772 1629
rect 3051 1611 3069 1665
rect 2592 1116 2610 1161
rect 2754 1116 2772 1161
rect 3051 1143 3069 1197
rect 4266 2727 4284 2772
rect 4428 2727 4446 2772
rect 4725 2754 4743 2808
rect 4266 2196 4284 2241
rect 4428 2196 4446 2241
rect 4725 2223 4743 2277
rect 5067 1593 5085 1638
rect 5229 1593 5247 1638
rect 5526 1620 5544 1674
rect 5067 1098 5085 1143
rect 5229 1098 5247 1143
rect 5526 1125 5544 1179
rect 2259 954 2277 1008
rect 2268 630 2286 684
rect 2592 675 2610 720
rect 2754 675 2772 720
rect 3051 702 3069 756
rect 5067 684 5085 729
rect 5229 684 5247 729
rect 5526 711 5544 765
rect 2592 261 2610 306
rect 2754 261 2772 306
rect 3051 288 3069 342
rect 3456 -216 3474 -171
rect 3618 -216 3636 -171
rect 3915 -189 3933 -135
rect 3456 -711 3474 -666
rect 3618 -711 3636 -666
rect 3915 -684 3933 -630
rect 3456 -1125 3474 -1080
rect 3618 -1125 3636 -1080
rect 3915 -1098 3933 -1044
rect 3456 -1656 3474 -1611
rect 3618 -1656 3636 -1611
rect 3915 -1629 3933 -1575
rect 3411 -2484 3429 -2439
rect 3573 -2484 3591 -2439
rect 3870 -2457 3888 -2403
rect 5067 153 5085 198
rect 5229 153 5247 198
rect 5526 180 5544 234
rect 6246 -171 6264 -126
rect 6408 -171 6426 -126
rect 6705 -144 6723 -90
rect 6246 -666 6264 -621
rect 6408 -666 6426 -621
rect 6705 -639 6723 -585
rect 6246 -1080 6264 -1035
rect 6408 -1080 6426 -1035
rect 6705 -1053 6723 -999
rect 5121 -2367 5139 -2322
rect 6246 -1611 6264 -1566
rect 6408 -1611 6426 -1566
rect 6705 -1584 6723 -1530
rect 5283 -2367 5301 -2322
rect 5580 -2340 5598 -2286
rect 5121 -2844 5139 -2799
rect 3411 -2979 3429 -2934
rect 3573 -2979 3591 -2934
rect 3870 -2952 3888 -2898
rect 5283 -2844 5301 -2799
rect 5580 -2817 5598 -2763
rect 5121 -3240 5139 -3195
rect 5283 -3240 5301 -3195
rect 5580 -3213 5598 -3159
rect 3411 -3393 3429 -3348
rect 3573 -3393 3591 -3348
rect 3870 -3366 3888 -3312
rect 5121 -3708 5139 -3663
rect 5283 -3708 5301 -3663
rect 5580 -3681 5598 -3627
rect 3411 -3924 3429 -3879
rect 3573 -3924 3591 -3879
rect 3870 -3897 3888 -3843
<< ndiffusion >>
rect 4680 6021 4725 6030
rect 4680 6003 4689 6021
rect 4716 6003 4725 6021
rect 4743 6003 4761 6030
rect 4788 6003 4797 6030
rect 4230 5967 4266 5976
rect 4230 5949 4239 5967
rect 4257 5949 4266 5967
rect 4284 5949 4428 5976
rect 4446 5958 4455 5976
rect 4473 5958 4482 5976
rect 4446 5949 4482 5958
rect 4680 5526 4725 5535
rect 4680 5508 4689 5526
rect 4716 5508 4725 5526
rect 4743 5508 4761 5535
rect 4788 5508 4797 5535
rect 4230 5472 4266 5481
rect 4230 5454 4239 5472
rect 4257 5454 4266 5472
rect 4284 5454 4428 5481
rect 4446 5463 4455 5481
rect 4473 5463 4482 5481
rect 4446 5454 4482 5463
rect 4680 5112 4725 5121
rect 4680 5094 4689 5112
rect 4716 5094 4725 5112
rect 4743 5094 4761 5121
rect 4788 5094 4797 5121
rect 4230 5058 4266 5067
rect 4230 5040 4239 5058
rect 4257 5040 4266 5058
rect 4284 5040 4428 5067
rect 4446 5049 4455 5067
rect 4473 5049 4482 5067
rect 4446 5040 4482 5049
rect 4680 4581 4725 4590
rect 4680 4563 4689 4581
rect 4716 4563 4725 4581
rect 4743 4563 4761 4590
rect 4788 4563 4797 4590
rect 4230 4527 4266 4536
rect 4230 4509 4239 4527
rect 4257 4509 4266 4527
rect 4284 4509 4428 4536
rect 4446 4518 4455 4536
rect 4473 4518 4482 4536
rect 4446 4509 4482 4518
rect 4680 3582 4725 3591
rect 4680 3564 4689 3582
rect 4716 3564 4725 3582
rect 4743 3564 4761 3591
rect 4788 3564 4797 3591
rect 4230 3528 4266 3537
rect 4230 3510 4239 3528
rect 4257 3510 4266 3528
rect 4284 3510 4428 3537
rect 4446 3519 4455 3537
rect 4473 3519 4482 3537
rect 4446 3510 4482 3519
rect 4680 3087 4725 3096
rect 4680 3069 4689 3087
rect 4716 3069 4725 3087
rect 4743 3069 4761 3096
rect 4788 3069 4797 3096
rect 4230 3033 4266 3042
rect 4230 3015 4239 3033
rect 4257 3015 4266 3033
rect 4284 3015 4428 3042
rect 4446 3024 4455 3042
rect 4473 3024 4482 3042
rect 4446 3015 4482 3024
rect 3663 2781 3672 2799
rect 3690 2781 3699 2799
rect 3663 2772 3699 2781
rect 3717 2781 3726 2799
rect 3717 2772 3744 2781
rect 3753 2781 3762 2799
rect 3780 2781 3789 2799
rect 3753 2772 3789 2781
rect 3807 2781 3816 2799
rect 3807 2772 3834 2781
rect 3879 2781 3888 2799
rect 3906 2781 3915 2799
rect 3879 2772 3915 2781
rect 3933 2781 3942 2799
rect 3960 2781 3969 2799
rect 3933 2772 3969 2781
rect 3006 1530 3051 1539
rect 3006 1512 3015 1530
rect 3042 1512 3051 1530
rect 3069 1512 3087 1539
rect 3114 1512 3123 1539
rect 2556 1476 2592 1485
rect 2556 1458 2565 1476
rect 2583 1458 2592 1476
rect 2610 1458 2754 1485
rect 2772 1467 2781 1485
rect 2799 1467 2808 1485
rect 2772 1458 2808 1467
rect 4680 2673 4725 2682
rect 4680 2655 4689 2673
rect 4716 2655 4725 2673
rect 4743 2655 4761 2682
rect 4788 2655 4797 2682
rect 4230 2619 4266 2628
rect 4230 2601 4239 2619
rect 4257 2601 4266 2619
rect 4284 2601 4428 2628
rect 4446 2610 4455 2628
rect 4473 2610 4482 2628
rect 4446 2601 4482 2610
rect 4680 2142 4725 2151
rect 4680 2124 4689 2142
rect 4716 2124 4725 2142
rect 4743 2124 4761 2151
rect 4788 2124 4797 2151
rect 4230 2088 4266 2097
rect 4230 2070 4239 2088
rect 4257 2070 4266 2088
rect 4284 2070 4428 2097
rect 4446 2079 4455 2097
rect 4473 2079 4482 2097
rect 4446 2070 4482 2079
rect 5481 1539 5526 1548
rect 5481 1521 5490 1539
rect 3006 1062 3051 1071
rect 3006 1044 3015 1062
rect 3042 1044 3051 1062
rect 3069 1044 3087 1071
rect 3114 1044 3123 1071
rect 5517 1521 5526 1539
rect 5544 1521 5562 1548
rect 5589 1521 5598 1548
rect 5031 1485 5067 1494
rect 5031 1467 5040 1485
rect 5058 1467 5067 1485
rect 5085 1467 5229 1494
rect 5247 1476 5256 1494
rect 5274 1476 5283 1494
rect 5247 1467 5283 1476
rect 5481 1044 5526 1053
rect 5481 1026 5490 1044
rect 2556 1008 2592 1017
rect 2556 990 2565 1008
rect 2583 990 2592 1008
rect 2610 990 2754 1017
rect 2772 999 2781 1017
rect 2799 999 2808 1017
rect 2772 990 2808 999
rect 2214 873 2259 882
rect 2214 855 2223 873
rect 2250 855 2259 873
rect 2277 855 2295 882
rect 2322 855 2331 882
rect 5517 1026 5526 1044
rect 5544 1026 5562 1053
rect 5589 1026 5598 1053
rect 5031 990 5067 999
rect 5031 972 5040 990
rect 5058 972 5067 990
rect 5085 972 5229 999
rect 5247 981 5256 999
rect 5274 981 5283 999
rect 5247 972 5283 981
rect 3006 621 3051 630
rect 3006 603 3015 621
rect 3042 603 3051 621
rect 3069 603 3087 630
rect 3114 603 3123 630
rect 2556 567 2592 576
rect 2223 549 2268 558
rect 2223 531 2232 549
rect 2259 531 2268 549
rect 2286 531 2304 558
rect 2331 531 2340 558
rect 2556 549 2565 567
rect 2583 549 2592 567
rect 2610 549 2727 576
rect 2745 549 2754 576
rect 2772 558 2781 576
rect 2799 558 2808 576
rect 2772 549 2808 558
rect 3006 207 3051 216
rect 3006 189 3015 207
rect 3042 189 3051 207
rect 3069 189 3087 216
rect 3114 189 3123 216
rect 2556 153 2592 162
rect 2556 135 2565 153
rect 2583 135 2592 153
rect 2610 135 2709 162
rect 2727 135 2754 162
rect 2772 144 2781 162
rect 2799 144 2808 162
rect 2772 135 2808 144
rect 3870 -270 3915 -261
rect 3870 -288 3879 -270
rect 3906 -288 3915 -270
rect 3933 -288 3951 -261
rect 3978 -288 3987 -261
rect 3420 -324 3456 -315
rect 3420 -342 3429 -324
rect 3447 -342 3456 -324
rect 3474 -342 3618 -315
rect 3636 -333 3645 -315
rect 3663 -333 3672 -315
rect 3636 -342 3672 -333
rect 3870 -765 3915 -756
rect 3870 -783 3879 -765
rect 3906 -783 3915 -765
rect 3933 -783 3951 -756
rect 3978 -783 3987 -756
rect 3420 -819 3456 -810
rect 3420 -837 3429 -819
rect 3447 -837 3456 -819
rect 3474 -837 3618 -810
rect 3636 -828 3645 -810
rect 3663 -828 3672 -810
rect 3636 -837 3672 -828
rect 3870 -1179 3915 -1170
rect 3870 -1197 3879 -1179
rect 3906 -1197 3915 -1179
rect 3933 -1197 3951 -1170
rect 3978 -1197 3987 -1170
rect 3420 -1233 3456 -1224
rect 3420 -1251 3429 -1233
rect 3447 -1251 3456 -1233
rect 3474 -1251 3618 -1224
rect 3636 -1242 3645 -1224
rect 3663 -1242 3672 -1224
rect 3636 -1251 3672 -1242
rect 3870 -1710 3915 -1701
rect 3870 -1728 3879 -1710
rect 3906 -1728 3915 -1710
rect 3933 -1728 3951 -1701
rect 3978 -1728 3987 -1701
rect 3420 -1764 3456 -1755
rect 3420 -1782 3429 -1764
rect 3447 -1782 3456 -1764
rect 3474 -1782 3618 -1755
rect 3636 -1773 3645 -1755
rect 3663 -1773 3672 -1755
rect 3636 -1782 3672 -1773
rect 3825 -2538 3870 -2529
rect 3825 -2556 3834 -2538
rect 3861 -2556 3870 -2538
rect 3888 -2556 3906 -2529
rect 3933 -2556 3942 -2529
rect 3375 -2592 3411 -2583
rect 3375 -2610 3384 -2592
rect 3402 -2610 3411 -2592
rect 3429 -2610 3573 -2583
rect 3591 -2601 3600 -2583
rect 3618 -2601 3627 -2583
rect 3591 -2610 3627 -2601
rect 5481 630 5526 639
rect 5481 612 5490 630
rect 5517 612 5526 630
rect 5544 612 5562 639
rect 5589 612 5598 639
rect 5031 576 5067 585
rect 5031 558 5040 576
rect 5058 558 5067 576
rect 5085 558 5229 585
rect 5247 567 5256 585
rect 5274 567 5283 585
rect 5247 558 5283 567
rect 5481 99 5526 108
rect 5481 81 5490 99
rect 5517 81 5526 99
rect 5544 81 5562 108
rect 5589 81 5598 108
rect 5031 45 5067 54
rect 5031 27 5040 45
rect 5058 27 5067 45
rect 5085 27 5229 54
rect 5247 36 5256 54
rect 5274 36 5283 54
rect 5247 27 5283 36
rect 6660 -225 6705 -216
rect 6660 -243 6669 -225
rect 6696 -243 6705 -225
rect 6723 -243 6741 -216
rect 6768 -243 6777 -216
rect 6210 -279 6246 -270
rect 6210 -297 6219 -279
rect 6237 -297 6246 -279
rect 6264 -297 6408 -270
rect 6426 -288 6435 -270
rect 6453 -288 6462 -270
rect 6426 -297 6462 -288
rect 6660 -720 6705 -711
rect 6660 -738 6669 -720
rect 6696 -738 6705 -720
rect 6723 -738 6741 -711
rect 6768 -738 6777 -711
rect 6210 -774 6246 -765
rect 6210 -792 6219 -774
rect 6237 -792 6246 -774
rect 6264 -792 6408 -765
rect 6426 -783 6435 -765
rect 6453 -783 6462 -765
rect 6426 -792 6462 -783
rect 6660 -1134 6705 -1125
rect 6660 -1152 6669 -1134
rect 6696 -1152 6705 -1134
rect 6723 -1152 6741 -1125
rect 6768 -1152 6777 -1125
rect 6210 -1188 6246 -1179
rect 6210 -1206 6219 -1188
rect 6237 -1206 6246 -1188
rect 6264 -1206 6408 -1179
rect 6426 -1197 6435 -1179
rect 6453 -1197 6462 -1179
rect 6426 -1206 6462 -1197
rect 6660 -1665 6705 -1656
rect 6660 -1683 6669 -1665
rect 6696 -1683 6705 -1665
rect 6723 -1683 6741 -1656
rect 6768 -1683 6777 -1656
rect 6210 -1719 6246 -1710
rect 6210 -1737 6219 -1719
rect 6237 -1737 6246 -1719
rect 6264 -1737 6408 -1710
rect 6426 -1728 6435 -1710
rect 6453 -1728 6462 -1710
rect 6426 -1737 6462 -1728
rect 5535 -2421 5580 -2412
rect 5535 -2439 5544 -2421
rect 5571 -2439 5580 -2421
rect 5598 -2439 5616 -2412
rect 5643 -2439 5652 -2412
rect 5085 -2475 5121 -2466
rect 5085 -2493 5094 -2475
rect 5112 -2493 5121 -2475
rect 5139 -2493 5283 -2466
rect 5301 -2484 5310 -2466
rect 5328 -2484 5337 -2466
rect 5301 -2493 5337 -2484
rect 5535 -2898 5580 -2889
rect 5535 -2916 5544 -2898
rect 5571 -2916 5580 -2898
rect 5598 -2916 5616 -2889
rect 5643 -2916 5652 -2889
rect 5085 -2952 5121 -2943
rect 5085 -2970 5094 -2952
rect 5112 -2970 5121 -2952
rect 5139 -2970 5283 -2943
rect 5301 -2961 5310 -2943
rect 5328 -2961 5337 -2943
rect 5301 -2970 5337 -2961
rect 3825 -3033 3870 -3024
rect 3825 -3051 3834 -3033
rect 3861 -3051 3870 -3033
rect 3888 -3051 3906 -3024
rect 3933 -3051 3942 -3024
rect 3375 -3087 3411 -3078
rect 3375 -3105 3384 -3087
rect 3402 -3105 3411 -3087
rect 3429 -3105 3573 -3078
rect 3591 -3096 3600 -3078
rect 3618 -3096 3627 -3078
rect 3591 -3105 3627 -3096
rect 5535 -3294 5580 -3285
rect 5535 -3312 5544 -3294
rect 5571 -3312 5580 -3294
rect 5598 -3312 5616 -3285
rect 5643 -3312 5652 -3285
rect 5085 -3348 5121 -3339
rect 5085 -3366 5094 -3348
rect 5112 -3366 5121 -3348
rect 5139 -3366 5283 -3339
rect 5301 -3357 5310 -3339
rect 5328 -3357 5337 -3339
rect 5301 -3366 5337 -3357
rect 3825 -3447 3870 -3438
rect 3825 -3465 3834 -3447
rect 3861 -3465 3870 -3447
rect 3888 -3465 3906 -3438
rect 3933 -3465 3942 -3438
rect 3375 -3501 3411 -3492
rect 3375 -3519 3384 -3501
rect 3402 -3519 3411 -3501
rect 3429 -3519 3573 -3492
rect 3591 -3510 3600 -3492
rect 3618 -3510 3627 -3492
rect 3591 -3519 3627 -3510
rect 5535 -3762 5580 -3753
rect 5535 -3780 5544 -3762
rect 5571 -3780 5580 -3762
rect 5598 -3780 5616 -3753
rect 5643 -3780 5652 -3753
rect 5085 -3816 5121 -3807
rect 5085 -3834 5094 -3816
rect 5112 -3834 5121 -3816
rect 5139 -3834 5283 -3807
rect 5301 -3825 5310 -3807
rect 5328 -3825 5337 -3807
rect 5301 -3834 5337 -3825
rect 3825 -3978 3870 -3969
rect 3825 -3996 3834 -3978
rect 3861 -3996 3870 -3978
rect 3888 -3996 3906 -3969
rect 3933 -3996 3942 -3969
rect 3375 -4032 3411 -4023
rect 3375 -4050 3384 -4032
rect 3402 -4050 3411 -4032
rect 3429 -4050 3573 -4023
rect 3591 -4041 3600 -4023
rect 3618 -4041 3627 -4023
rect 3591 -4050 3627 -4041
<< pdiffusion >>
rect 4680 6129 4689 6156
rect 4716 6129 4725 6156
rect 4230 6111 4266 6120
rect 4230 6093 4239 6111
rect 4257 6093 4266 6111
rect 4230 6075 4266 6093
rect 4284 6102 4347 6120
rect 4284 6084 4293 6102
rect 4311 6084 4347 6102
rect 4284 6075 4347 6084
rect 4383 6111 4428 6120
rect 4383 6093 4392 6111
rect 4410 6093 4428 6111
rect 4383 6075 4428 6093
rect 4446 6111 4482 6120
rect 4446 6093 4455 6111
rect 4473 6093 4482 6111
rect 4680 6102 4725 6129
rect 4743 6147 4797 6156
rect 4743 6120 4761 6147
rect 4788 6120 4797 6147
rect 4743 6102 4797 6120
rect 4446 6075 4482 6093
rect 4680 5634 4689 5661
rect 4716 5634 4725 5661
rect 4230 5616 4266 5625
rect 4230 5598 4239 5616
rect 4257 5598 4266 5616
rect 4230 5580 4266 5598
rect 4284 5607 4347 5625
rect 4284 5589 4293 5607
rect 4311 5589 4347 5607
rect 4284 5580 4347 5589
rect 4383 5616 4428 5625
rect 4383 5598 4392 5616
rect 4410 5598 4428 5616
rect 4383 5580 4428 5598
rect 4446 5616 4482 5625
rect 4446 5598 4455 5616
rect 4473 5598 4482 5616
rect 4680 5607 4725 5634
rect 4743 5652 4797 5661
rect 4743 5625 4761 5652
rect 4788 5625 4797 5652
rect 4743 5607 4797 5625
rect 4446 5580 4482 5598
rect 4680 5220 4689 5247
rect 4716 5220 4725 5247
rect 4230 5202 4266 5211
rect 4230 5184 4239 5202
rect 4257 5184 4266 5202
rect 4230 5166 4266 5184
rect 4284 5193 4347 5211
rect 4284 5175 4293 5193
rect 4311 5175 4347 5193
rect 4284 5166 4347 5175
rect 4383 5202 4428 5211
rect 4383 5184 4392 5202
rect 4410 5184 4428 5202
rect 4383 5166 4428 5184
rect 4446 5202 4482 5211
rect 4446 5184 4455 5202
rect 4473 5184 4482 5202
rect 4680 5193 4725 5220
rect 4743 5238 4797 5247
rect 4743 5211 4761 5238
rect 4788 5211 4797 5238
rect 4743 5193 4797 5211
rect 4446 5166 4482 5184
rect 4680 4689 4689 4716
rect 4716 4689 4725 4716
rect 4230 4671 4266 4680
rect 4230 4653 4239 4671
rect 4257 4653 4266 4671
rect 4230 4635 4266 4653
rect 4284 4662 4347 4680
rect 4284 4644 4293 4662
rect 4311 4644 4347 4662
rect 4284 4635 4347 4644
rect 4383 4671 4428 4680
rect 4383 4653 4392 4671
rect 4410 4653 4428 4671
rect 4383 4635 4428 4653
rect 4446 4671 4482 4680
rect 4446 4653 4455 4671
rect 4473 4653 4482 4671
rect 4680 4662 4725 4689
rect 4743 4707 4797 4716
rect 4743 4680 4761 4707
rect 4788 4680 4797 4707
rect 4743 4662 4797 4680
rect 4446 4635 4482 4653
rect 4680 3690 4689 3717
rect 4716 3690 4725 3717
rect 4230 3672 4266 3681
rect 4230 3654 4239 3672
rect 4257 3654 4266 3672
rect 4230 3636 4266 3654
rect 4284 3663 4347 3681
rect 4284 3645 4293 3663
rect 4311 3645 4347 3663
rect 4284 3636 4347 3645
rect 4383 3672 4428 3681
rect 4383 3654 4392 3672
rect 4410 3654 4428 3672
rect 4383 3636 4428 3654
rect 4446 3672 4482 3681
rect 4446 3654 4455 3672
rect 4473 3654 4482 3672
rect 4680 3663 4725 3690
rect 4743 3708 4797 3717
rect 4743 3681 4761 3708
rect 4788 3681 4797 3708
rect 4743 3663 4797 3681
rect 4446 3636 4482 3654
rect 4680 3195 4689 3222
rect 4716 3195 4725 3222
rect 4230 3177 4266 3186
rect 4230 3159 4239 3177
rect 4257 3159 4266 3177
rect 4230 3141 4266 3159
rect 4284 3168 4347 3186
rect 4284 3150 4293 3168
rect 4311 3150 4347 3168
rect 4284 3141 4347 3150
rect 4383 3177 4428 3186
rect 4383 3159 4392 3177
rect 4410 3159 4428 3177
rect 4383 3141 4428 3159
rect 4446 3177 4482 3186
rect 4446 3159 4455 3177
rect 4473 3159 4482 3177
rect 4680 3168 4725 3195
rect 4743 3213 4797 3222
rect 4743 3186 4761 3213
rect 4788 3186 4797 3213
rect 4743 3168 4797 3186
rect 4446 3141 4482 3159
rect 3654 2925 3699 2934
rect 3654 2907 3663 2925
rect 3681 2907 3699 2925
rect 3654 2889 3699 2907
rect 3717 2889 3789 2934
rect 3807 2916 3834 2934
rect 3807 2898 3816 2916
rect 3807 2889 3834 2898
rect 3879 2925 3915 2934
rect 3879 2907 3888 2925
rect 3906 2907 3915 2925
rect 3879 2889 3915 2907
rect 3933 2916 3969 2934
rect 3933 2898 3942 2916
rect 3960 2898 3969 2916
rect 3933 2889 3969 2898
rect 3006 1638 3015 1665
rect 3042 1638 3051 1665
rect 2556 1620 2592 1629
rect 2556 1602 2565 1620
rect 2583 1602 2592 1620
rect 2556 1584 2592 1602
rect 2610 1611 2673 1629
rect 2610 1593 2619 1611
rect 2637 1593 2673 1611
rect 2610 1584 2673 1593
rect 2709 1620 2754 1629
rect 2709 1602 2718 1620
rect 2736 1602 2754 1620
rect 2709 1584 2754 1602
rect 2772 1620 2808 1629
rect 2772 1602 2781 1620
rect 2799 1602 2808 1620
rect 3006 1611 3051 1638
rect 3069 1656 3123 1665
rect 3069 1629 3087 1656
rect 3114 1629 3123 1656
rect 3069 1611 3123 1629
rect 2772 1584 2808 1602
rect 3006 1170 3015 1197
rect 3042 1170 3051 1197
rect 2556 1152 2592 1161
rect 2556 1134 2565 1152
rect 2583 1134 2592 1152
rect 2556 1116 2592 1134
rect 2610 1143 2673 1161
rect 2610 1125 2619 1143
rect 2637 1125 2673 1143
rect 2610 1116 2673 1125
rect 2709 1152 2754 1161
rect 2709 1134 2718 1152
rect 2736 1134 2754 1152
rect 2709 1116 2754 1134
rect 2772 1152 2808 1161
rect 2772 1134 2781 1152
rect 2799 1134 2808 1152
rect 3006 1143 3051 1170
rect 3069 1188 3123 1197
rect 3069 1161 3087 1188
rect 3114 1161 3123 1188
rect 3069 1143 3123 1161
rect 2772 1116 2808 1134
rect 4680 2781 4689 2808
rect 4716 2781 4725 2808
rect 4230 2763 4266 2772
rect 4230 2745 4239 2763
rect 4257 2745 4266 2763
rect 4230 2727 4266 2745
rect 4284 2754 4347 2772
rect 4284 2736 4293 2754
rect 4311 2736 4347 2754
rect 4284 2727 4347 2736
rect 4383 2763 4428 2772
rect 4383 2745 4392 2763
rect 4410 2745 4428 2763
rect 4383 2727 4428 2745
rect 4446 2763 4482 2772
rect 4446 2745 4455 2763
rect 4473 2745 4482 2763
rect 4680 2754 4725 2781
rect 4743 2799 4797 2808
rect 4743 2772 4761 2799
rect 4788 2772 4797 2799
rect 4743 2754 4797 2772
rect 4446 2727 4482 2745
rect 4680 2250 4689 2277
rect 4716 2250 4725 2277
rect 4230 2232 4266 2241
rect 4230 2214 4239 2232
rect 4257 2214 4266 2232
rect 4230 2196 4266 2214
rect 4284 2223 4347 2241
rect 4284 2205 4293 2223
rect 4311 2205 4347 2223
rect 4284 2196 4347 2205
rect 4383 2232 4428 2241
rect 4383 2214 4392 2232
rect 4410 2214 4428 2232
rect 4383 2196 4428 2214
rect 4446 2232 4482 2241
rect 4446 2214 4455 2232
rect 4473 2214 4482 2232
rect 4680 2223 4725 2250
rect 4743 2268 4797 2277
rect 4743 2241 4761 2268
rect 4788 2241 4797 2268
rect 4743 2223 4797 2241
rect 4446 2196 4482 2214
rect 5481 1647 5490 1674
rect 5517 1647 5526 1674
rect 5031 1629 5067 1638
rect 5031 1611 5040 1629
rect 5058 1611 5067 1629
rect 5031 1593 5067 1611
rect 5085 1620 5148 1638
rect 5085 1602 5094 1620
rect 5112 1602 5148 1620
rect 5085 1593 5148 1602
rect 5184 1629 5229 1638
rect 5184 1611 5193 1629
rect 5211 1611 5229 1629
rect 5184 1593 5229 1611
rect 5247 1629 5283 1638
rect 5247 1611 5256 1629
rect 5274 1611 5283 1629
rect 5481 1620 5526 1647
rect 5544 1665 5598 1674
rect 5544 1638 5562 1665
rect 5589 1638 5598 1665
rect 5544 1620 5598 1638
rect 5247 1593 5283 1611
rect 5481 1152 5490 1179
rect 5517 1152 5526 1179
rect 5031 1134 5067 1143
rect 5031 1116 5040 1134
rect 5058 1116 5067 1134
rect 5031 1098 5067 1116
rect 5085 1125 5148 1143
rect 5085 1107 5094 1125
rect 5112 1107 5148 1125
rect 5085 1098 5148 1107
rect 5184 1134 5229 1143
rect 5184 1116 5193 1134
rect 5211 1116 5229 1134
rect 5184 1098 5229 1116
rect 5247 1134 5283 1143
rect 5247 1116 5256 1134
rect 5274 1116 5283 1134
rect 5481 1125 5526 1152
rect 5544 1170 5598 1179
rect 5544 1143 5562 1170
rect 5589 1143 5598 1170
rect 5544 1125 5598 1143
rect 5247 1098 5283 1116
rect 2214 981 2223 1008
rect 2250 981 2259 1008
rect 2214 954 2259 981
rect 2277 999 2331 1008
rect 2277 972 2295 999
rect 2322 972 2331 999
rect 2277 954 2331 972
rect 3006 729 3015 756
rect 3042 729 3051 756
rect 2556 711 2592 720
rect 2556 693 2565 711
rect 2583 693 2592 711
rect 2223 657 2232 684
rect 2259 657 2268 684
rect 2223 630 2268 657
rect 2286 675 2340 684
rect 2556 675 2592 693
rect 2610 702 2673 720
rect 2610 684 2619 702
rect 2637 684 2673 702
rect 2610 675 2673 684
rect 2709 711 2754 720
rect 2709 693 2718 711
rect 2736 693 2754 711
rect 2709 675 2754 693
rect 2772 711 2808 720
rect 2772 693 2781 711
rect 2799 693 2808 711
rect 3006 702 3051 729
rect 3069 747 3123 756
rect 3069 720 3087 747
rect 3114 720 3123 747
rect 3069 702 3123 720
rect 2772 675 2808 693
rect 2286 648 2304 675
rect 2331 648 2340 675
rect 2286 630 2340 648
rect 5481 738 5490 765
rect 5517 738 5526 765
rect 5031 720 5067 729
rect 5031 702 5040 720
rect 5058 702 5067 720
rect 5031 684 5067 702
rect 5085 711 5148 729
rect 5085 693 5094 711
rect 5112 693 5148 711
rect 5085 684 5148 693
rect 5184 720 5229 729
rect 5184 702 5193 720
rect 5211 702 5229 720
rect 5184 684 5229 702
rect 5247 720 5283 729
rect 5247 702 5256 720
rect 5274 702 5283 720
rect 5481 711 5526 738
rect 5544 756 5598 765
rect 5544 729 5562 756
rect 5589 729 5598 756
rect 5544 711 5598 729
rect 5247 684 5283 702
rect 3006 315 3015 342
rect 3042 315 3051 342
rect 2556 297 2592 306
rect 2556 279 2565 297
rect 2583 279 2592 297
rect 2556 261 2592 279
rect 2610 288 2673 306
rect 2610 270 2619 288
rect 2637 270 2673 288
rect 2610 261 2673 270
rect 2709 297 2754 306
rect 2709 279 2718 297
rect 2736 279 2754 297
rect 2709 261 2754 279
rect 2772 297 2808 306
rect 2772 279 2781 297
rect 2799 279 2808 297
rect 3006 288 3051 315
rect 3069 333 3123 342
rect 3069 306 3087 333
rect 3114 306 3123 333
rect 3069 288 3123 306
rect 2772 261 2808 279
rect 3870 -162 3879 -135
rect 3906 -162 3915 -135
rect 3420 -180 3456 -171
rect 3420 -198 3429 -180
rect 3447 -198 3456 -180
rect 3420 -216 3456 -198
rect 3474 -189 3537 -171
rect 3474 -207 3483 -189
rect 3501 -207 3537 -189
rect 3474 -216 3537 -207
rect 3573 -180 3618 -171
rect 3573 -198 3582 -180
rect 3600 -198 3618 -180
rect 3573 -216 3618 -198
rect 3636 -180 3672 -171
rect 3636 -198 3645 -180
rect 3663 -198 3672 -180
rect 3870 -189 3915 -162
rect 3933 -144 3987 -135
rect 3933 -171 3951 -144
rect 3978 -171 3987 -144
rect 3933 -189 3987 -171
rect 3636 -216 3672 -198
rect 3870 -657 3879 -630
rect 3906 -657 3915 -630
rect 3420 -675 3456 -666
rect 3420 -693 3429 -675
rect 3447 -693 3456 -675
rect 3420 -711 3456 -693
rect 3474 -684 3537 -666
rect 3474 -702 3483 -684
rect 3501 -702 3537 -684
rect 3474 -711 3537 -702
rect 3573 -675 3618 -666
rect 3573 -693 3582 -675
rect 3600 -693 3618 -675
rect 3573 -711 3618 -693
rect 3636 -675 3672 -666
rect 3636 -693 3645 -675
rect 3663 -693 3672 -675
rect 3870 -684 3915 -657
rect 3933 -639 3987 -630
rect 3933 -666 3951 -639
rect 3978 -666 3987 -639
rect 3933 -684 3987 -666
rect 3636 -711 3672 -693
rect 3870 -1071 3879 -1044
rect 3906 -1071 3915 -1044
rect 3420 -1089 3456 -1080
rect 3420 -1107 3429 -1089
rect 3447 -1107 3456 -1089
rect 3420 -1125 3456 -1107
rect 3474 -1098 3537 -1080
rect 3474 -1116 3483 -1098
rect 3501 -1116 3537 -1098
rect 3474 -1125 3537 -1116
rect 3573 -1089 3618 -1080
rect 3573 -1107 3582 -1089
rect 3600 -1107 3618 -1089
rect 3573 -1125 3618 -1107
rect 3636 -1089 3672 -1080
rect 3636 -1107 3645 -1089
rect 3663 -1107 3672 -1089
rect 3870 -1098 3915 -1071
rect 3933 -1053 3987 -1044
rect 3933 -1080 3951 -1053
rect 3978 -1080 3987 -1053
rect 3933 -1098 3987 -1080
rect 3636 -1125 3672 -1107
rect 3870 -1602 3879 -1575
rect 3906 -1602 3915 -1575
rect 3420 -1620 3456 -1611
rect 3420 -1638 3429 -1620
rect 3447 -1638 3456 -1620
rect 3420 -1656 3456 -1638
rect 3474 -1629 3537 -1611
rect 3474 -1647 3483 -1629
rect 3501 -1647 3537 -1629
rect 3474 -1656 3537 -1647
rect 3573 -1620 3618 -1611
rect 3573 -1638 3582 -1620
rect 3600 -1638 3618 -1620
rect 3573 -1656 3618 -1638
rect 3636 -1620 3672 -1611
rect 3636 -1638 3645 -1620
rect 3663 -1638 3672 -1620
rect 3870 -1629 3915 -1602
rect 3933 -1584 3987 -1575
rect 3933 -1611 3951 -1584
rect 3978 -1611 3987 -1584
rect 3933 -1629 3987 -1611
rect 3636 -1656 3672 -1638
rect 3825 -2430 3834 -2403
rect 3861 -2430 3870 -2403
rect 3375 -2448 3411 -2439
rect 3375 -2466 3384 -2448
rect 3402 -2466 3411 -2448
rect 3375 -2484 3411 -2466
rect 3429 -2457 3492 -2439
rect 3429 -2475 3438 -2457
rect 3456 -2475 3492 -2457
rect 3429 -2484 3492 -2475
rect 3528 -2448 3573 -2439
rect 3528 -2466 3537 -2448
rect 3555 -2466 3573 -2448
rect 3528 -2484 3573 -2466
rect 3591 -2448 3627 -2439
rect 3591 -2466 3600 -2448
rect 3618 -2466 3627 -2448
rect 3825 -2457 3870 -2430
rect 3888 -2412 3942 -2403
rect 3888 -2439 3906 -2412
rect 3933 -2439 3942 -2412
rect 3888 -2457 3942 -2439
rect 3591 -2484 3627 -2466
rect 5481 207 5490 234
rect 5517 207 5526 234
rect 5031 189 5067 198
rect 5031 171 5040 189
rect 5058 171 5067 189
rect 5031 153 5067 171
rect 5085 180 5148 198
rect 5085 162 5094 180
rect 5112 162 5148 180
rect 5085 153 5148 162
rect 5184 189 5229 198
rect 5184 171 5193 189
rect 5211 171 5229 189
rect 5184 153 5229 171
rect 5247 189 5283 198
rect 5247 171 5256 189
rect 5274 171 5283 189
rect 5481 180 5526 207
rect 5544 225 5598 234
rect 5544 198 5562 225
rect 5589 198 5598 225
rect 5544 180 5598 198
rect 5247 153 5283 171
rect 6660 -117 6669 -90
rect 6696 -117 6705 -90
rect 6210 -135 6246 -126
rect 6210 -153 6219 -135
rect 6237 -153 6246 -135
rect 6210 -171 6246 -153
rect 6264 -144 6327 -126
rect 6264 -162 6273 -144
rect 6291 -162 6327 -144
rect 6264 -171 6327 -162
rect 6363 -135 6408 -126
rect 6363 -153 6372 -135
rect 6390 -153 6408 -135
rect 6363 -171 6408 -153
rect 6426 -135 6462 -126
rect 6426 -153 6435 -135
rect 6453 -153 6462 -135
rect 6660 -144 6705 -117
rect 6723 -99 6777 -90
rect 6723 -126 6741 -99
rect 6768 -126 6777 -99
rect 6723 -144 6777 -126
rect 6426 -171 6462 -153
rect 6660 -612 6669 -585
rect 6696 -612 6705 -585
rect 6210 -630 6246 -621
rect 6210 -648 6219 -630
rect 6237 -648 6246 -630
rect 6210 -666 6246 -648
rect 6264 -639 6327 -621
rect 6264 -657 6273 -639
rect 6291 -657 6327 -639
rect 6264 -666 6327 -657
rect 6363 -630 6408 -621
rect 6363 -648 6372 -630
rect 6390 -648 6408 -630
rect 6363 -666 6408 -648
rect 6426 -630 6462 -621
rect 6426 -648 6435 -630
rect 6453 -648 6462 -630
rect 6660 -639 6705 -612
rect 6723 -594 6777 -585
rect 6723 -621 6741 -594
rect 6768 -621 6777 -594
rect 6723 -639 6777 -621
rect 6426 -666 6462 -648
rect 6660 -1026 6669 -999
rect 6696 -1026 6705 -999
rect 6210 -1044 6246 -1035
rect 6210 -1062 6219 -1044
rect 6237 -1062 6246 -1044
rect 6210 -1080 6246 -1062
rect 6264 -1053 6327 -1035
rect 6264 -1071 6273 -1053
rect 6291 -1071 6327 -1053
rect 6264 -1080 6327 -1071
rect 6363 -1044 6408 -1035
rect 6363 -1062 6372 -1044
rect 6390 -1062 6408 -1044
rect 6363 -1080 6408 -1062
rect 6426 -1044 6462 -1035
rect 6426 -1062 6435 -1044
rect 6453 -1062 6462 -1044
rect 6660 -1053 6705 -1026
rect 6723 -1008 6777 -999
rect 6723 -1035 6741 -1008
rect 6768 -1035 6777 -1008
rect 6723 -1053 6777 -1035
rect 6426 -1080 6462 -1062
rect 5085 -2331 5121 -2322
rect 5085 -2349 5094 -2331
rect 5112 -2349 5121 -2331
rect 5085 -2367 5121 -2349
rect 5139 -2340 5202 -2322
rect 5139 -2358 5148 -2340
rect 5166 -2358 5202 -2340
rect 5139 -2367 5202 -2358
rect 6660 -1557 6669 -1530
rect 6696 -1557 6705 -1530
rect 6210 -1575 6246 -1566
rect 6210 -1593 6219 -1575
rect 6237 -1593 6246 -1575
rect 6210 -1611 6246 -1593
rect 6264 -1584 6327 -1566
rect 6264 -1602 6273 -1584
rect 6291 -1602 6327 -1584
rect 6264 -1611 6327 -1602
rect 6363 -1575 6408 -1566
rect 6363 -1593 6372 -1575
rect 6390 -1593 6408 -1575
rect 6363 -1611 6408 -1593
rect 6426 -1575 6462 -1566
rect 6426 -1593 6435 -1575
rect 6453 -1593 6462 -1575
rect 6660 -1584 6705 -1557
rect 6723 -1539 6777 -1530
rect 6723 -1566 6741 -1539
rect 6768 -1566 6777 -1539
rect 6723 -1584 6777 -1566
rect 6426 -1611 6462 -1593
rect 5535 -2313 5544 -2286
rect 5571 -2313 5580 -2286
rect 5238 -2331 5283 -2322
rect 5238 -2349 5247 -2331
rect 5265 -2349 5283 -2331
rect 5238 -2367 5283 -2349
rect 5301 -2331 5337 -2322
rect 5301 -2349 5310 -2331
rect 5328 -2349 5337 -2331
rect 5535 -2340 5580 -2313
rect 5598 -2295 5652 -2286
rect 5598 -2322 5616 -2295
rect 5643 -2322 5652 -2295
rect 5598 -2340 5652 -2322
rect 5301 -2367 5337 -2349
rect 5085 -2808 5121 -2799
rect 5085 -2826 5094 -2808
rect 5112 -2826 5121 -2808
rect 5085 -2844 5121 -2826
rect 5139 -2817 5202 -2799
rect 5139 -2835 5148 -2817
rect 5166 -2835 5202 -2817
rect 5139 -2844 5202 -2835
rect 3825 -2925 3834 -2898
rect 3861 -2925 3870 -2898
rect 3375 -2943 3411 -2934
rect 3375 -2961 3384 -2943
rect 3402 -2961 3411 -2943
rect 3375 -2979 3411 -2961
rect 3429 -2952 3492 -2934
rect 3429 -2970 3438 -2952
rect 3456 -2970 3492 -2952
rect 3429 -2979 3492 -2970
rect 3528 -2943 3573 -2934
rect 3528 -2961 3537 -2943
rect 3555 -2961 3573 -2943
rect 3528 -2979 3573 -2961
rect 3591 -2943 3627 -2934
rect 3591 -2961 3600 -2943
rect 3618 -2961 3627 -2943
rect 3825 -2952 3870 -2925
rect 3888 -2907 3942 -2898
rect 3888 -2934 3906 -2907
rect 3933 -2934 3942 -2907
rect 3888 -2952 3942 -2934
rect 3591 -2979 3627 -2961
rect 5535 -2790 5544 -2763
rect 5571 -2790 5580 -2763
rect 5238 -2808 5283 -2799
rect 5238 -2826 5247 -2808
rect 5265 -2826 5283 -2808
rect 5238 -2844 5283 -2826
rect 5301 -2808 5337 -2799
rect 5301 -2826 5310 -2808
rect 5328 -2826 5337 -2808
rect 5535 -2817 5580 -2790
rect 5598 -2772 5652 -2763
rect 5598 -2799 5616 -2772
rect 5643 -2799 5652 -2772
rect 5598 -2817 5652 -2799
rect 5301 -2844 5337 -2826
rect 5535 -3186 5544 -3159
rect 5571 -3186 5580 -3159
rect 5085 -3204 5121 -3195
rect 5085 -3222 5094 -3204
rect 5112 -3222 5121 -3204
rect 5085 -3240 5121 -3222
rect 5139 -3213 5202 -3195
rect 5139 -3231 5148 -3213
rect 5166 -3231 5202 -3213
rect 5139 -3240 5202 -3231
rect 5238 -3204 5283 -3195
rect 5238 -3222 5247 -3204
rect 5265 -3222 5283 -3204
rect 5238 -3240 5283 -3222
rect 5301 -3204 5337 -3195
rect 5301 -3222 5310 -3204
rect 5328 -3222 5337 -3204
rect 5535 -3213 5580 -3186
rect 5598 -3168 5652 -3159
rect 5598 -3195 5616 -3168
rect 5643 -3195 5652 -3168
rect 5598 -3213 5652 -3195
rect 5301 -3240 5337 -3222
rect 3825 -3339 3834 -3312
rect 3861 -3339 3870 -3312
rect 3375 -3357 3411 -3348
rect 3375 -3375 3384 -3357
rect 3402 -3375 3411 -3357
rect 3375 -3393 3411 -3375
rect 3429 -3366 3492 -3348
rect 3429 -3384 3438 -3366
rect 3456 -3384 3492 -3366
rect 3429 -3393 3492 -3384
rect 3528 -3357 3573 -3348
rect 3528 -3375 3537 -3357
rect 3555 -3375 3573 -3357
rect 3528 -3393 3573 -3375
rect 3591 -3357 3627 -3348
rect 3591 -3375 3600 -3357
rect 3618 -3375 3627 -3357
rect 3825 -3366 3870 -3339
rect 3888 -3321 3942 -3312
rect 3888 -3348 3906 -3321
rect 3933 -3348 3942 -3321
rect 3888 -3366 3942 -3348
rect 3591 -3393 3627 -3375
rect 5535 -3654 5544 -3627
rect 5571 -3654 5580 -3627
rect 5085 -3672 5121 -3663
rect 5085 -3690 5094 -3672
rect 5112 -3690 5121 -3672
rect 5085 -3708 5121 -3690
rect 5139 -3681 5202 -3663
rect 5139 -3699 5148 -3681
rect 5166 -3699 5202 -3681
rect 5139 -3708 5202 -3699
rect 5238 -3672 5283 -3663
rect 5238 -3690 5247 -3672
rect 5265 -3690 5283 -3672
rect 5238 -3708 5283 -3690
rect 5301 -3672 5337 -3663
rect 5301 -3690 5310 -3672
rect 5328 -3690 5337 -3672
rect 5535 -3681 5580 -3654
rect 5598 -3636 5652 -3627
rect 5598 -3663 5616 -3636
rect 5643 -3663 5652 -3636
rect 5598 -3681 5652 -3663
rect 5301 -3708 5337 -3690
rect 3825 -3870 3834 -3843
rect 3861 -3870 3870 -3843
rect 3375 -3888 3411 -3879
rect 3375 -3906 3384 -3888
rect 3402 -3906 3411 -3888
rect 3375 -3924 3411 -3906
rect 3429 -3897 3492 -3879
rect 3429 -3915 3438 -3897
rect 3456 -3915 3492 -3897
rect 3429 -3924 3492 -3915
rect 3528 -3888 3573 -3879
rect 3528 -3906 3537 -3888
rect 3555 -3906 3573 -3888
rect 3528 -3924 3573 -3906
rect 3591 -3888 3627 -3879
rect 3591 -3906 3600 -3888
rect 3618 -3906 3627 -3888
rect 3825 -3897 3870 -3870
rect 3888 -3852 3942 -3843
rect 3888 -3879 3906 -3852
rect 3933 -3879 3942 -3852
rect 3888 -3897 3942 -3879
rect 3591 -3924 3627 -3906
<< ndcontact >>
rect 4689 5994 4716 6021
rect 4761 6003 4788 6030
rect 4239 5949 4257 5967
rect 4455 5958 4473 5976
rect 4689 5499 4716 5526
rect 4761 5508 4788 5535
rect 4239 5454 4257 5472
rect 4455 5463 4473 5481
rect 4689 5085 4716 5112
rect 4761 5094 4788 5121
rect 4239 5040 4257 5058
rect 4455 5049 4473 5067
rect 4689 4554 4716 4581
rect 4761 4563 4788 4590
rect 4239 4509 4257 4527
rect 4455 4518 4473 4536
rect 4689 3555 4716 3582
rect 4761 3564 4788 3591
rect 4239 3510 4257 3528
rect 4455 3519 4473 3537
rect 4689 3060 4716 3087
rect 4761 3069 4788 3096
rect 4239 3015 4257 3033
rect 4455 3024 4473 3042
rect 3672 2781 3690 2799
rect 3726 2781 3744 2799
rect 3762 2781 3780 2799
rect 3816 2781 3834 2799
rect 3888 2781 3906 2799
rect 3942 2781 3960 2799
rect 3015 1503 3042 1530
rect 3087 1512 3114 1539
rect 2565 1458 2583 1476
rect 2781 1467 2799 1485
rect 4689 2646 4716 2673
rect 4761 2655 4788 2682
rect 4239 2601 4257 2619
rect 4455 2610 4473 2628
rect 4689 2115 4716 2142
rect 4761 2124 4788 2151
rect 4239 2070 4257 2088
rect 4455 2079 4473 2097
rect 3015 1035 3042 1062
rect 3087 1044 3114 1071
rect 5490 1512 5517 1539
rect 5562 1521 5589 1548
rect 5040 1467 5058 1485
rect 5256 1476 5274 1494
rect 2565 990 2583 1008
rect 2781 999 2799 1017
rect 2223 846 2250 873
rect 2295 855 2322 882
rect 5490 1017 5517 1044
rect 5562 1026 5589 1053
rect 5040 972 5058 990
rect 5256 981 5274 999
rect 3015 594 3042 621
rect 3087 603 3114 630
rect 2232 522 2259 549
rect 2304 531 2331 558
rect 2565 549 2583 567
rect 2781 558 2799 576
rect 3015 180 3042 207
rect 3087 189 3114 216
rect 2565 135 2583 153
rect 2781 144 2799 162
rect 3879 -297 3906 -270
rect 3951 -288 3978 -261
rect 3429 -342 3447 -324
rect 3645 -333 3663 -315
rect 3879 -792 3906 -765
rect 3951 -783 3978 -756
rect 3429 -837 3447 -819
rect 3645 -828 3663 -810
rect 3879 -1206 3906 -1179
rect 3951 -1197 3978 -1170
rect 3429 -1251 3447 -1233
rect 3645 -1242 3663 -1224
rect 3879 -1737 3906 -1710
rect 3951 -1728 3978 -1701
rect 3429 -1782 3447 -1764
rect 3645 -1773 3663 -1755
rect 3834 -2565 3861 -2538
rect 3906 -2556 3933 -2529
rect 3384 -2610 3402 -2592
rect 3600 -2601 3618 -2583
rect 5490 603 5517 630
rect 5562 612 5589 639
rect 5040 558 5058 576
rect 5256 567 5274 585
rect 5490 72 5517 99
rect 5562 81 5589 108
rect 5040 27 5058 45
rect 5256 36 5274 54
rect 6669 -252 6696 -225
rect 6741 -243 6768 -216
rect 6219 -297 6237 -279
rect 6435 -288 6453 -270
rect 6669 -747 6696 -720
rect 6741 -738 6768 -711
rect 6219 -792 6237 -774
rect 6435 -783 6453 -765
rect 6669 -1161 6696 -1134
rect 6741 -1152 6768 -1125
rect 6219 -1206 6237 -1188
rect 6435 -1197 6453 -1179
rect 6669 -1692 6696 -1665
rect 6741 -1683 6768 -1656
rect 6219 -1737 6237 -1719
rect 6435 -1728 6453 -1710
rect 5544 -2448 5571 -2421
rect 5616 -2439 5643 -2412
rect 5094 -2493 5112 -2475
rect 5310 -2484 5328 -2466
rect 5544 -2925 5571 -2898
rect 5616 -2916 5643 -2889
rect 5094 -2970 5112 -2952
rect 5310 -2961 5328 -2943
rect 3834 -3060 3861 -3033
rect 3906 -3051 3933 -3024
rect 3384 -3105 3402 -3087
rect 3600 -3096 3618 -3078
rect 5544 -3321 5571 -3294
rect 5616 -3312 5643 -3285
rect 5094 -3366 5112 -3348
rect 5310 -3357 5328 -3339
rect 3834 -3474 3861 -3447
rect 3906 -3465 3933 -3438
rect 3384 -3519 3402 -3501
rect 3600 -3510 3618 -3492
rect 5544 -3789 5571 -3762
rect 5616 -3780 5643 -3753
rect 5094 -3834 5112 -3816
rect 5310 -3825 5328 -3807
rect 3834 -4005 3861 -3978
rect 3906 -3996 3933 -3969
rect 3384 -4050 3402 -4032
rect 3600 -4041 3618 -4023
<< pdcontact >>
rect 4689 6129 4716 6156
rect 4239 6093 4257 6111
rect 4293 6084 4311 6102
rect 4392 6093 4410 6111
rect 4455 6093 4473 6111
rect 4761 6120 4788 6147
rect 4689 5634 4716 5661
rect 4239 5598 4257 5616
rect 4293 5589 4311 5607
rect 4392 5598 4410 5616
rect 4455 5598 4473 5616
rect 4761 5625 4788 5652
rect 4689 5220 4716 5247
rect 4239 5184 4257 5202
rect 4293 5175 4311 5193
rect 4392 5184 4410 5202
rect 4455 5184 4473 5202
rect 4761 5211 4788 5238
rect 4689 4689 4716 4716
rect 4239 4653 4257 4671
rect 4293 4644 4311 4662
rect 4392 4653 4410 4671
rect 4455 4653 4473 4671
rect 4761 4680 4788 4707
rect 4689 3690 4716 3717
rect 4239 3654 4257 3672
rect 4293 3645 4311 3663
rect 4392 3654 4410 3672
rect 4455 3654 4473 3672
rect 4761 3681 4788 3708
rect 4689 3195 4716 3222
rect 4239 3159 4257 3177
rect 4293 3150 4311 3168
rect 4392 3159 4410 3177
rect 4455 3159 4473 3177
rect 4761 3186 4788 3213
rect 3663 2907 3681 2925
rect 3816 2898 3834 2916
rect 3888 2907 3906 2925
rect 3942 2898 3960 2916
rect 3015 1638 3042 1665
rect 2565 1602 2583 1620
rect 2619 1593 2637 1611
rect 2718 1602 2736 1620
rect 2781 1602 2799 1620
rect 3087 1629 3114 1656
rect 3015 1170 3042 1197
rect 2565 1134 2583 1152
rect 2619 1125 2637 1143
rect 2718 1134 2736 1152
rect 2781 1134 2799 1152
rect 3087 1161 3114 1188
rect 4689 2781 4716 2808
rect 4239 2745 4257 2763
rect 4293 2736 4311 2754
rect 4392 2745 4410 2763
rect 4455 2745 4473 2763
rect 4761 2772 4788 2799
rect 4689 2250 4716 2277
rect 4239 2214 4257 2232
rect 4293 2205 4311 2223
rect 4392 2214 4410 2232
rect 4455 2214 4473 2232
rect 4761 2241 4788 2268
rect 5490 1647 5517 1674
rect 5040 1611 5058 1629
rect 5094 1602 5112 1620
rect 5193 1611 5211 1629
rect 5256 1611 5274 1629
rect 5562 1638 5589 1665
rect 5490 1152 5517 1179
rect 5040 1116 5058 1134
rect 5094 1107 5112 1125
rect 5193 1116 5211 1134
rect 5256 1116 5274 1134
rect 5562 1143 5589 1170
rect 2223 981 2250 1008
rect 2295 972 2322 999
rect 3015 729 3042 756
rect 2565 693 2583 711
rect 2232 657 2259 684
rect 2619 684 2637 702
rect 2718 693 2736 711
rect 2781 693 2799 711
rect 3087 720 3114 747
rect 2304 648 2331 675
rect 5490 738 5517 765
rect 5040 702 5058 720
rect 5094 693 5112 711
rect 5193 702 5211 720
rect 5256 702 5274 720
rect 5562 729 5589 756
rect 3015 315 3042 342
rect 2565 279 2583 297
rect 2619 270 2637 288
rect 2718 279 2736 297
rect 2781 279 2799 297
rect 3087 306 3114 333
rect 3879 -162 3906 -135
rect 3429 -198 3447 -180
rect 3483 -207 3501 -189
rect 3582 -198 3600 -180
rect 3645 -198 3663 -180
rect 3951 -171 3978 -144
rect 3879 -657 3906 -630
rect 3429 -693 3447 -675
rect 3483 -702 3501 -684
rect 3582 -693 3600 -675
rect 3645 -693 3663 -675
rect 3951 -666 3978 -639
rect 3879 -1071 3906 -1044
rect 3429 -1107 3447 -1089
rect 3483 -1116 3501 -1098
rect 3582 -1107 3600 -1089
rect 3645 -1107 3663 -1089
rect 3951 -1080 3978 -1053
rect 3879 -1602 3906 -1575
rect 3429 -1638 3447 -1620
rect 3483 -1647 3501 -1629
rect 3582 -1638 3600 -1620
rect 3645 -1638 3663 -1620
rect 3951 -1611 3978 -1584
rect 3834 -2430 3861 -2403
rect 3384 -2466 3402 -2448
rect 3438 -2475 3456 -2457
rect 3537 -2466 3555 -2448
rect 3600 -2466 3618 -2448
rect 3906 -2439 3933 -2412
rect 5490 207 5517 234
rect 5040 171 5058 189
rect 5094 162 5112 180
rect 5193 171 5211 189
rect 5256 171 5274 189
rect 5562 198 5589 225
rect 6669 -117 6696 -90
rect 6219 -153 6237 -135
rect 6273 -162 6291 -144
rect 6372 -153 6390 -135
rect 6435 -153 6453 -135
rect 6741 -126 6768 -99
rect 6669 -612 6696 -585
rect 6219 -648 6237 -630
rect 6273 -657 6291 -639
rect 6372 -648 6390 -630
rect 6435 -648 6453 -630
rect 6741 -621 6768 -594
rect 6669 -1026 6696 -999
rect 6219 -1062 6237 -1044
rect 6273 -1071 6291 -1053
rect 6372 -1062 6390 -1044
rect 6435 -1062 6453 -1044
rect 6741 -1035 6768 -1008
rect 5094 -2349 5112 -2331
rect 5148 -2358 5166 -2340
rect 6669 -1557 6696 -1530
rect 6219 -1593 6237 -1575
rect 6273 -1602 6291 -1584
rect 6372 -1593 6390 -1575
rect 6435 -1593 6453 -1575
rect 6741 -1566 6768 -1539
rect 5544 -2313 5571 -2286
rect 5247 -2349 5265 -2331
rect 5310 -2349 5328 -2331
rect 5616 -2322 5643 -2295
rect 5094 -2826 5112 -2808
rect 5148 -2835 5166 -2817
rect 3834 -2925 3861 -2898
rect 3384 -2961 3402 -2943
rect 3438 -2970 3456 -2952
rect 3537 -2961 3555 -2943
rect 3600 -2961 3618 -2943
rect 3906 -2934 3933 -2907
rect 5544 -2790 5571 -2763
rect 5247 -2826 5265 -2808
rect 5310 -2826 5328 -2808
rect 5616 -2799 5643 -2772
rect 5544 -3186 5571 -3159
rect 5094 -3222 5112 -3204
rect 5148 -3231 5166 -3213
rect 5247 -3222 5265 -3204
rect 5310 -3222 5328 -3204
rect 5616 -3195 5643 -3168
rect 3834 -3339 3861 -3312
rect 3384 -3375 3402 -3357
rect 3438 -3384 3456 -3366
rect 3537 -3375 3555 -3357
rect 3600 -3375 3618 -3357
rect 3906 -3348 3933 -3321
rect 5544 -3654 5571 -3627
rect 5094 -3690 5112 -3672
rect 5148 -3699 5166 -3681
rect 5247 -3690 5265 -3672
rect 5310 -3690 5328 -3672
rect 5616 -3663 5643 -3636
rect 3834 -3870 3861 -3843
rect 3384 -3906 3402 -3888
rect 3438 -3915 3456 -3897
rect 3537 -3906 3555 -3888
rect 3600 -3906 3618 -3888
rect 3906 -3879 3933 -3852
<< polysilicon >>
rect 4725 6156 4743 6273
rect 4266 6120 4284 6147
rect 4428 6120 4446 6147
rect 4266 6012 4284 6075
rect 4095 5994 4284 6012
rect 4428 6003 4446 6075
rect 4725 6066 4743 6102
rect 4734 6039 4743 6066
rect 4725 6030 4743 6039
rect 4095 5517 4113 5994
rect 4266 5976 4284 5994
rect 4725 5985 4743 6003
rect 4428 5976 4446 5985
rect 4266 5940 4284 5949
rect 4428 5940 4446 5949
rect 4725 5661 4743 5778
rect 4266 5625 4284 5652
rect 4428 5625 4446 5652
rect 4266 5517 4284 5580
rect 4095 5499 4284 5517
rect 4428 5508 4446 5580
rect 4725 5571 4743 5607
rect 4734 5544 4743 5571
rect 4725 5535 4743 5544
rect 4095 5283 4113 5499
rect 4266 5481 4284 5499
rect 4725 5490 4743 5508
rect 4428 5481 4446 5490
rect 4266 5445 4284 5454
rect 4428 5445 4446 5454
rect 4068 5265 4113 5283
rect 4095 5094 4113 5265
rect 4725 5247 4743 5364
rect 4266 5211 4284 5238
rect 4428 5211 4446 5238
rect 4266 5094 4284 5166
rect 4428 5094 4446 5166
rect 4725 5157 4743 5193
rect 4734 5130 4743 5157
rect 4725 5121 4743 5130
rect 4095 5076 4284 5094
rect 4725 5076 4743 5094
rect 4095 4572 4113 5076
rect 4266 5067 4284 5076
rect 4428 5067 4446 5076
rect 4266 5031 4284 5040
rect 4428 5031 4446 5040
rect 4725 4716 4743 4833
rect 4266 4680 4284 4707
rect 4428 4680 4446 4707
rect 4266 4572 4284 4635
rect 4095 4554 4284 4572
rect 4428 4563 4446 4635
rect 4725 4626 4743 4662
rect 4734 4599 4743 4626
rect 4725 4590 4743 4599
rect 4095 3573 4113 4554
rect 4266 4536 4284 4554
rect 4725 4545 4743 4563
rect 4428 4536 4446 4545
rect 4266 4500 4284 4509
rect 4428 4500 4446 4509
rect 4725 3717 4743 3834
rect 4266 3681 4284 3708
rect 4428 3681 4446 3708
rect 4266 3573 4284 3636
rect 4095 3555 4284 3573
rect 4428 3564 4446 3636
rect 4725 3627 4743 3663
rect 4734 3600 4743 3627
rect 4725 3591 4743 3600
rect 4095 3078 4113 3555
rect 4266 3537 4284 3555
rect 4725 3546 4743 3564
rect 4428 3537 4446 3546
rect 4266 3501 4284 3510
rect 4428 3501 4446 3510
rect 4725 3222 4743 3339
rect 4266 3186 4284 3213
rect 4428 3186 4446 3213
rect 4266 3078 4284 3141
rect 4095 3060 4284 3078
rect 4428 3069 4446 3141
rect 4725 3132 4743 3168
rect 4734 3105 4743 3132
rect 4725 3096 4743 3105
rect 3699 2934 3717 2952
rect 3789 2934 3807 2952
rect 3915 2934 3933 2952
rect 3699 2844 3717 2889
rect 3465 2817 3717 2844
rect 3051 1665 3069 1782
rect 2592 1629 2610 1656
rect 2754 1629 2772 1656
rect 2592 1530 2610 1584
rect 2754 1512 2772 1584
rect 3051 1575 3069 1611
rect 3465 1584 3492 2817
rect 3699 2799 3717 2817
rect 3789 2799 3807 2889
rect 3915 2844 3933 2889
rect 4095 2844 4113 3060
rect 4266 3042 4284 3060
rect 4725 3051 4743 3069
rect 4428 3042 4446 3051
rect 4266 3006 4284 3015
rect 4428 3006 4446 3015
rect 3924 2826 3933 2844
rect 4005 2826 4113 2844
rect 3915 2799 3933 2826
rect 3699 2763 3717 2772
rect 3060 1548 3069 1575
rect 3159 1557 3492 1584
rect 3051 1539 3069 1548
rect 2592 1485 2610 1512
rect 3051 1494 3069 1512
rect 2754 1485 2772 1494
rect 2592 1449 2610 1458
rect 2754 1449 2772 1458
rect 2124 1197 2520 1215
rect 3051 1197 3069 1314
rect 2124 918 2142 1197
rect 2502 1053 2520 1197
rect 2592 1161 2610 1188
rect 2754 1161 2772 1188
rect 2592 1053 2610 1116
rect 2502 1035 2610 1053
rect 2259 1008 2277 1026
rect 2592 1017 2610 1035
rect 2754 1044 2772 1116
rect 3051 1107 3069 1143
rect 3789 1116 3807 2772
rect 3915 2763 3933 2772
rect 4095 2655 4113 2826
rect 4725 2808 4743 2925
rect 4266 2772 4284 2799
rect 4428 2772 4446 2799
rect 4266 2655 4284 2727
rect 4428 2655 4446 2727
rect 4725 2718 4743 2754
rect 4734 2691 4743 2718
rect 4725 2682 4743 2691
rect 4095 2637 4284 2655
rect 4725 2637 4743 2655
rect 4095 2133 4113 2637
rect 4266 2628 4284 2637
rect 4428 2628 4446 2637
rect 4266 2592 4284 2601
rect 4428 2592 4446 2601
rect 4725 2277 4743 2394
rect 4266 2241 4284 2268
rect 4428 2241 4446 2268
rect 4266 2133 4284 2196
rect 4095 2115 4284 2133
rect 4428 2124 4446 2196
rect 4725 2187 4743 2223
rect 4734 2160 4743 2187
rect 4725 2151 4743 2160
rect 4266 2097 4284 2115
rect 4725 2106 4743 2124
rect 4428 2097 4446 2106
rect 4266 2061 4284 2070
rect 4428 2061 4446 2070
rect 5526 1674 5544 1791
rect 5067 1638 5085 1665
rect 5229 1638 5247 1665
rect 5067 1530 5085 1593
rect 3060 1080 3069 1107
rect 3159 1089 3807 1116
rect 4896 1512 5085 1530
rect 5229 1521 5247 1593
rect 5526 1584 5544 1620
rect 5535 1557 5544 1584
rect 5526 1548 5544 1557
rect 3051 1071 3069 1080
rect 3051 1026 3069 1044
rect 4896 1035 4914 1512
rect 5067 1494 5085 1512
rect 5526 1503 5544 1521
rect 5229 1494 5247 1503
rect 5067 1458 5085 1467
rect 5229 1458 5247 1467
rect 5526 1179 5544 1296
rect 5067 1143 5085 1170
rect 5229 1143 5247 1170
rect 5067 1035 5085 1098
rect 2754 1017 2772 1026
rect 4896 1017 5085 1035
rect 5229 1026 5247 1098
rect 5526 1089 5544 1125
rect 5535 1062 5544 1089
rect 5526 1053 5544 1062
rect 2592 981 2610 990
rect 2754 981 2772 990
rect 2259 918 2277 954
rect 2007 891 2277 918
rect 2007 54 2025 891
rect 2259 882 2277 891
rect 2259 837 2277 855
rect 3051 756 3069 873
rect 2592 720 2610 747
rect 2754 720 2772 747
rect 2268 684 2286 702
rect 2592 630 2610 675
rect 2268 594 2286 630
rect 2061 567 2286 594
rect 2592 576 2610 612
rect 2754 603 2772 675
rect 3051 666 3069 702
rect 4896 675 4914 1017
rect 5067 999 5085 1017
rect 5526 1008 5544 1026
rect 5229 999 5247 1008
rect 5067 963 5085 972
rect 5229 963 5247 972
rect 5526 765 5544 882
rect 5067 729 5085 756
rect 5229 729 5247 756
rect 3060 639 3069 666
rect 3150 648 4914 675
rect 3051 630 3069 639
rect 2727 585 2772 603
rect 3051 585 3069 603
rect 2727 576 2745 585
rect 2754 576 2772 585
rect 2061 450 2079 567
rect 2268 558 2286 567
rect 2592 540 2610 549
rect 2268 513 2286 531
rect 2727 450 2745 549
rect 2754 540 2772 549
rect 2061 432 2745 450
rect 2448 225 2466 432
rect 3051 342 3069 459
rect 2592 306 2610 333
rect 2754 306 2772 333
rect 2592 225 2610 261
rect 2448 207 2610 225
rect 2592 162 2610 207
rect 2754 189 2772 261
rect 3051 252 3069 288
rect 3060 225 3069 252
rect 3132 234 3303 261
rect 3051 216 3069 225
rect 2709 171 2772 189
rect 3051 171 3069 189
rect 2709 162 2727 171
rect 2754 162 2772 171
rect 2592 126 2610 135
rect 2709 54 2727 135
rect 2754 126 2772 135
rect 2007 36 2727 54
rect 3285 -279 3303 234
rect 3915 -135 3933 -18
rect 3456 -171 3474 -144
rect 3618 -171 3636 -144
rect 3456 -279 3474 -216
rect 3285 -297 3474 -279
rect 3618 -288 3636 -216
rect 3915 -225 3933 -189
rect 3924 -252 3933 -225
rect 4005 -243 4617 -216
rect 3915 -261 3933 -252
rect 3285 -774 3303 -297
rect 3456 -315 3474 -297
rect 3915 -306 3933 -288
rect 3618 -315 3636 -306
rect 3456 -351 3474 -342
rect 3618 -351 3636 -342
rect 3915 -630 3933 -513
rect 3456 -666 3474 -639
rect 3618 -666 3636 -639
rect 3456 -774 3474 -711
rect 3285 -792 3474 -774
rect 3618 -783 3636 -711
rect 3915 -720 3933 -684
rect 3924 -747 3933 -720
rect 3915 -756 3933 -747
rect 3285 -1197 3303 -792
rect 3456 -810 3474 -792
rect 3915 -801 3933 -783
rect 3618 -810 3636 -801
rect 3456 -846 3474 -837
rect 3618 -846 3636 -837
rect 3915 -1044 3933 -927
rect 3456 -1080 3474 -1053
rect 3618 -1080 3636 -1053
rect 3456 -1197 3474 -1125
rect 3618 -1197 3636 -1125
rect 3915 -1134 3933 -1098
rect 3924 -1161 3933 -1134
rect 3915 -1170 3933 -1161
rect 3285 -1215 3474 -1197
rect 3915 -1215 3933 -1197
rect 3285 -1683 3303 -1215
rect 3456 -1224 3474 -1215
rect 3618 -1224 3636 -1215
rect 3456 -1260 3474 -1251
rect 3618 -1260 3636 -1251
rect 3915 -1575 3933 -1458
rect 3456 -1611 3474 -1584
rect 3618 -1611 3636 -1584
rect 3240 -1701 3303 -1683
rect 3240 -2547 3258 -1701
rect 3285 -1719 3303 -1701
rect 3456 -1719 3474 -1656
rect 3285 -1737 3474 -1719
rect 3618 -1728 3636 -1656
rect 3915 -1665 3933 -1629
rect 3924 -1692 3933 -1665
rect 3915 -1701 3933 -1692
rect 3456 -1755 3474 -1737
rect 3915 -1746 3933 -1728
rect 3618 -1755 3636 -1746
rect 3456 -1791 3474 -1782
rect 3618 -1791 3636 -1782
rect 4014 -2142 4032 -1530
rect 4383 -2223 4401 -576
rect 3636 -2241 4401 -2223
rect 3870 -2403 3888 -2286
rect 3411 -2439 3429 -2412
rect 3573 -2439 3591 -2412
rect 3411 -2547 3429 -2484
rect 3240 -2565 3429 -2547
rect 3240 -3042 3258 -2565
rect 3411 -2583 3429 -2565
rect 3573 -2556 3591 -2484
rect 3870 -2493 3888 -2457
rect 3879 -2520 3888 -2493
rect 3960 -2502 4320 -2484
rect 3870 -2529 3888 -2520
rect 3870 -2574 3888 -2556
rect 3573 -2583 3591 -2574
rect 3411 -2619 3429 -2610
rect 3573 -2619 3591 -2610
rect 4473 -2691 4491 -963
rect 4599 -1341 4617 -243
rect 4806 -729 4824 648
rect 4896 612 4914 648
rect 5067 612 5085 684
rect 5229 612 5247 684
rect 5526 675 5544 711
rect 5535 648 5544 675
rect 5526 639 5544 648
rect 4896 594 5085 612
rect 5526 594 5544 612
rect 4896 90 4914 594
rect 5067 585 5085 594
rect 5229 585 5247 594
rect 5067 549 5085 558
rect 5229 549 5247 558
rect 5526 234 5544 351
rect 5067 198 5085 225
rect 5229 198 5247 225
rect 5067 90 5085 153
rect 4896 72 5085 90
rect 5229 81 5247 153
rect 5526 144 5544 180
rect 5535 117 5544 144
rect 5526 108 5544 117
rect 5067 54 5085 72
rect 5526 63 5544 81
rect 5229 54 5247 63
rect 5067 18 5085 27
rect 5229 18 5247 27
rect 6705 -90 6723 27
rect 6246 -126 6264 -99
rect 6408 -126 6426 -99
rect 6246 -234 6264 -171
rect 6075 -252 6264 -234
rect 6408 -243 6426 -171
rect 6705 -180 6723 -144
rect 6714 -207 6723 -180
rect 6705 -216 6723 -207
rect 5211 -378 5940 -360
rect 5211 -549 5229 -378
rect 6075 -729 6093 -252
rect 6246 -270 6264 -252
rect 6705 -261 6723 -243
rect 6408 -270 6426 -261
rect 6246 -306 6264 -297
rect 6408 -306 6426 -297
rect 6705 -585 6723 -468
rect 6246 -621 6264 -594
rect 6408 -621 6426 -594
rect 6246 -729 6264 -666
rect 4806 -747 6264 -729
rect 6408 -738 6426 -666
rect 6705 -675 6723 -639
rect 6714 -702 6723 -675
rect 6705 -711 6723 -702
rect 5067 -954 5913 -936
rect 6075 -1152 6093 -747
rect 6246 -765 6264 -747
rect 6705 -756 6723 -738
rect 6408 -765 6426 -756
rect 6246 -801 6264 -792
rect 6408 -801 6426 -792
rect 6705 -999 6723 -882
rect 6246 -1035 6264 -1008
rect 6408 -1035 6426 -1008
rect 6246 -1152 6264 -1080
rect 6408 -1152 6426 -1080
rect 6705 -1089 6723 -1053
rect 6714 -1116 6723 -1089
rect 6705 -1125 6723 -1116
rect 6075 -1170 6264 -1152
rect 6705 -1170 6723 -1152
rect 4599 -1359 5229 -1341
rect 4671 -2655 4689 -1971
rect 5121 -2322 5139 -2295
rect 5121 -2412 5139 -2367
rect 4851 -2430 5139 -2412
rect 4851 -2484 4869 -2430
rect 5121 -2466 5139 -2430
rect 5211 -2439 5229 -1359
rect 6075 -1674 6093 -1170
rect 6246 -1179 6264 -1170
rect 6408 -1179 6426 -1170
rect 6246 -1215 6264 -1206
rect 6408 -1215 6426 -1206
rect 6705 -1530 6723 -1413
rect 6246 -1566 6264 -1539
rect 6408 -1566 6426 -1539
rect 6246 -1674 6264 -1611
rect 6075 -1692 6264 -1674
rect 6408 -1683 6426 -1611
rect 6705 -1620 6723 -1584
rect 6714 -1647 6723 -1620
rect 6705 -1656 6723 -1647
rect 6246 -1710 6264 -1692
rect 6705 -1701 6723 -1683
rect 6408 -1710 6426 -1701
rect 6246 -1746 6264 -1737
rect 6408 -1746 6426 -1737
rect 5580 -2286 5598 -2169
rect 5283 -2322 5301 -2295
rect 5283 -2439 5301 -2367
rect 5580 -2376 5598 -2340
rect 5589 -2403 5598 -2376
rect 5580 -2412 5598 -2403
rect 5211 -2457 5301 -2439
rect 5580 -2457 5598 -2439
rect 5283 -2466 5301 -2457
rect 5121 -2502 5139 -2493
rect 5283 -2502 5301 -2493
rect 4671 -2673 5229 -2655
rect 3582 -2709 4491 -2691
rect 3870 -2898 3888 -2781
rect 5121 -2799 5139 -2772
rect 5121 -2898 5139 -2844
rect 3411 -2934 3429 -2907
rect 3573 -2934 3591 -2907
rect 4167 -2916 5139 -2898
rect 3411 -3042 3429 -2979
rect 3240 -3060 3429 -3042
rect 3573 -3051 3591 -2979
rect 3870 -2988 3888 -2952
rect 4167 -2979 4185 -2916
rect 5121 -2943 5139 -2916
rect 5211 -2916 5229 -2673
rect 5580 -2763 5598 -2646
rect 5283 -2799 5301 -2772
rect 5283 -2916 5301 -2844
rect 5580 -2853 5598 -2817
rect 5589 -2880 5598 -2853
rect 5580 -2889 5598 -2880
rect 5211 -2934 5301 -2916
rect 5580 -2934 5598 -2916
rect 5283 -2943 5301 -2934
rect 5121 -2979 5139 -2970
rect 5283 -2979 5301 -2970
rect 3879 -3015 3888 -2988
rect 3960 -3006 4185 -2979
rect 3870 -3024 3888 -3015
rect 3240 -3465 3258 -3060
rect 3411 -3078 3429 -3060
rect 3870 -3069 3888 -3051
rect 3573 -3078 3591 -3069
rect 3411 -3114 3429 -3105
rect 3573 -3114 3591 -3105
rect 5580 -3159 5598 -3042
rect 5121 -3195 5139 -3168
rect 5283 -3195 5301 -3168
rect 3870 -3312 3888 -3195
rect 5121 -3294 5139 -3240
rect 4230 -3312 5085 -3294
rect 3411 -3348 3429 -3321
rect 3573 -3348 3591 -3321
rect 3411 -3465 3429 -3393
rect 3573 -3465 3591 -3393
rect 3870 -3402 3888 -3366
rect 4230 -3393 4248 -3312
rect 5121 -3339 5139 -3312
rect 5283 -3312 5301 -3240
rect 5580 -3249 5598 -3213
rect 5589 -3276 5598 -3249
rect 5580 -3285 5598 -3276
rect 5580 -3330 5598 -3312
rect 5283 -3339 5301 -3330
rect 5121 -3375 5139 -3366
rect 5283 -3375 5301 -3366
rect 3879 -3429 3888 -3402
rect 3960 -3420 4248 -3393
rect 3870 -3438 3888 -3429
rect 3240 -3483 3429 -3465
rect 3870 -3483 3888 -3465
rect 3240 -3987 3258 -3483
rect 3411 -3492 3429 -3483
rect 3573 -3492 3591 -3483
rect 3411 -3528 3429 -3519
rect 3573 -3528 3591 -3519
rect 5580 -3627 5598 -3510
rect 5121 -3663 5139 -3636
rect 5283 -3663 5301 -3636
rect 3870 -3843 3888 -3726
rect 5121 -3762 5139 -3708
rect 5112 -3780 5139 -3762
rect 5121 -3807 5139 -3780
rect 5283 -3780 5301 -3708
rect 5580 -3717 5598 -3681
rect 5589 -3744 5598 -3717
rect 5580 -3753 5598 -3744
rect 5580 -3798 5598 -3780
rect 5283 -3807 5301 -3798
rect 5121 -3843 5139 -3834
rect 5283 -3843 5301 -3834
rect 3411 -3879 3429 -3852
rect 3573 -3879 3591 -3852
rect 3411 -3987 3429 -3924
rect 3240 -4005 3429 -3987
rect 3573 -3996 3591 -3924
rect 3870 -3933 3888 -3897
rect 3879 -3960 3888 -3933
rect 3870 -3969 3888 -3960
rect 3411 -4023 3429 -4005
rect 3870 -4014 3888 -3996
rect 3573 -4023 3591 -4014
rect 3411 -4059 3429 -4050
rect 3573 -4059 3591 -4050
<< polycontact >>
rect 4707 6039 4734 6066
rect 4419 5985 4446 6003
rect 4707 5544 4734 5571
rect 4419 5490 4446 5508
rect 4707 5130 4734 5157
rect 4419 5076 4446 5094
rect 4707 4599 4734 4626
rect 4419 4545 4446 4563
rect 4707 3600 4734 3627
rect 4419 3546 4446 3564
rect 4707 3105 4734 3132
rect 2583 1512 2610 1530
rect 4419 3051 4446 3069
rect 3915 2826 3924 2844
rect 3960 2826 4005 2844
rect 3033 1548 3060 1575
rect 3114 1557 3159 1584
rect 2736 1494 2772 1512
rect 4707 2691 4734 2718
rect 4419 2637 4446 2655
rect 4707 2160 4734 2187
rect 4419 2106 4446 2124
rect 3033 1080 3060 1107
rect 3123 1089 3159 1116
rect 5508 1557 5535 1584
rect 2754 1026 2772 1044
rect 5220 1503 5247 1521
rect 5508 1062 5535 1089
rect 2592 612 2610 630
rect 5220 1008 5247 1026
rect 3033 639 3060 666
rect 3114 648 3150 675
rect 3033 225 3060 252
rect 3096 234 3132 261
rect 3897 -252 3924 -225
rect 3978 -243 4005 -216
rect 3609 -306 3636 -288
rect 4383 -576 4401 -549
rect 3897 -747 3924 -720
rect 3600 -801 3636 -783
rect 3897 -1161 3924 -1134
rect 3591 -1215 3636 -1197
rect 4014 -1530 4032 -1503
rect 3897 -1692 3924 -1665
rect 3591 -1746 3636 -1728
rect 4014 -2169 4032 -2142
rect 3564 -2241 3636 -2223
rect 4473 -963 4491 -936
rect 3852 -2520 3879 -2493
rect 3933 -2502 3960 -2484
rect 4320 -2502 4365 -2484
rect 3573 -2574 3591 -2556
rect 5508 648 5535 675
rect 5220 594 5247 612
rect 5508 117 5535 144
rect 5220 63 5247 81
rect 6687 -207 6714 -180
rect 5940 -378 5967 -360
rect 5211 -567 5229 -549
rect 6399 -261 6426 -243
rect 6687 -702 6714 -675
rect 5022 -954 5067 -936
rect 5913 -954 5931 -936
rect 6399 -756 6426 -738
rect 6687 -1116 6714 -1089
rect 6399 -1170 6426 -1152
rect 4671 -1971 4689 -1935
rect 6687 -1647 6714 -1620
rect 6399 -1701 6426 -1683
rect 5562 -2403 5589 -2376
rect 4851 -2502 4869 -2484
rect 3528 -2709 3582 -2691
rect 5562 -2880 5589 -2853
rect 3852 -3015 3879 -2988
rect 3924 -3006 3960 -2979
rect 3555 -3069 3591 -3051
rect 5085 -3312 5139 -3294
rect 5562 -3276 5589 -3249
rect 5283 -3330 5301 -3312
rect 3852 -3429 3879 -3402
rect 3933 -3420 3960 -3393
rect 3564 -3483 3591 -3465
rect 5067 -3780 5112 -3762
rect 5562 -3744 5589 -3717
rect 5283 -3798 5301 -3780
rect 3852 -3960 3879 -3933
rect 3564 -4014 3591 -3996
<< metal1 >>
rect 4689 6210 4923 6228
rect 4689 6183 4716 6210
rect 4068 6165 4716 6183
rect 4239 6111 4257 6165
rect 4392 6111 4410 6165
rect 4689 6156 4716 6165
rect 4293 6030 4311 6084
rect 4455 6030 4473 6093
rect 4761 6075 4788 6120
rect 4617 6039 4707 6066
rect 4761 6048 4815 6075
rect 4617 6030 4635 6039
rect 4293 6012 4635 6030
rect 4761 6030 4788 6048
rect 4410 5985 4419 6003
rect 4455 5976 4473 6012
rect 4689 5967 4716 5994
rect 4239 5931 4257 5949
rect 4689 5949 4788 5967
rect 4689 5931 4725 5949
rect 4131 5913 4725 5931
rect 4131 5436 4149 5913
rect 4905 5733 4923 6210
rect 4689 5715 4923 5733
rect 4689 5688 4716 5715
rect 4239 5670 4716 5688
rect 4239 5616 4257 5670
rect 4392 5616 4410 5670
rect 4689 5661 4716 5670
rect 4293 5535 4311 5589
rect 4455 5535 4473 5598
rect 4761 5580 4788 5625
rect 4617 5544 4707 5571
rect 4761 5553 4815 5580
rect 4617 5535 4635 5544
rect 4293 5517 4635 5535
rect 4761 5535 4788 5553
rect 4410 5490 4419 5508
rect 4455 5481 4473 5517
rect 4689 5472 4716 5499
rect 4239 5436 4257 5454
rect 4689 5454 4788 5472
rect 4689 5436 4725 5454
rect 4131 5418 4725 5436
rect 4131 5193 4149 5418
rect 4905 5319 4923 5715
rect 4689 5301 4923 5319
rect 4689 5274 4716 5301
rect 4068 5175 4149 5193
rect 4239 5256 4716 5274
rect 4239 5202 4257 5256
rect 4392 5202 4410 5256
rect 4689 5247 4716 5256
rect 4131 5022 4149 5175
rect 4293 5121 4311 5175
rect 4455 5121 4473 5184
rect 4761 5166 4788 5211
rect 4617 5130 4707 5157
rect 4761 5139 4815 5166
rect 4617 5121 4635 5130
rect 4293 5103 4635 5121
rect 4761 5121 4788 5139
rect 4410 5076 4419 5094
rect 4455 5067 4473 5103
rect 4689 5058 4716 5085
rect 4239 5022 4257 5040
rect 4689 5040 4788 5058
rect 4689 5022 4725 5040
rect 4131 5004 4725 5022
rect -315 4878 378 4896
rect 4131 4536 4149 5004
rect 4905 4788 4923 5301
rect 4689 4770 4923 4788
rect 4689 4743 4716 4770
rect 4239 4725 4716 4743
rect 4239 4671 4257 4725
rect 4392 4671 4410 4725
rect 4689 4716 4716 4725
rect 4293 4590 4311 4644
rect 4455 4590 4473 4653
rect 4761 4635 4788 4680
rect 4617 4599 4707 4626
rect 4761 4608 4815 4635
rect 4617 4590 4635 4599
rect 4293 4572 4635 4590
rect 4761 4590 4788 4608
rect 4410 4545 4419 4563
rect 4455 4536 4473 4572
rect 4689 4527 4716 4554
rect 4239 4491 4257 4509
rect 4689 4509 4788 4527
rect 4689 4491 4725 4509
rect 4149 4473 4725 4491
rect -216 4338 -45 4356
rect 4905 3789 4923 4770
rect 4689 3771 4923 3789
rect 4689 3744 4716 3771
rect 3888 3726 4716 3744
rect 3888 3582 3906 3726
rect 4239 3672 4257 3726
rect 4392 3672 4410 3726
rect 4689 3717 4716 3726
rect 2997 3564 3906 3582
rect 4293 3591 4311 3645
rect 4455 3591 4473 3654
rect 4761 3636 4788 3681
rect 4617 3600 4707 3627
rect 4761 3609 4815 3636
rect 4617 3591 4635 3600
rect 4293 3573 4635 3591
rect 4761 3591 4788 3609
rect 2997 1854 3015 3564
rect 3888 2979 3906 3564
rect 4455 3537 4473 3573
rect 4689 3528 4716 3555
rect 4239 3492 4257 3510
rect 4689 3510 4788 3528
rect 4689 3492 4725 3510
rect 4149 3474 4725 3492
rect 4131 2997 4149 3402
rect 4905 3294 4923 3771
rect 4689 3276 4923 3294
rect 4689 3249 4716 3276
rect 4239 3231 4716 3249
rect 4239 3177 4257 3231
rect 4392 3177 4410 3231
rect 4689 3222 4716 3231
rect 4293 3096 4311 3150
rect 4455 3096 4473 3159
rect 4761 3141 4788 3186
rect 4617 3105 4707 3132
rect 4761 3114 4815 3141
rect 4617 3096 4635 3105
rect 4293 3078 4635 3096
rect 4761 3096 4788 3114
rect 4410 3051 4419 3069
rect 4455 3042 4473 3078
rect 4689 3033 4716 3060
rect 4239 2997 4257 3015
rect 4689 3015 4788 3033
rect 4689 2997 4725 3015
rect 4131 2979 4725 2997
rect 3663 2961 3933 2979
rect 3663 2925 3681 2961
rect 3888 2925 3906 2961
rect 3816 2844 3834 2898
rect 3726 2826 3915 2844
rect 3726 2799 3744 2826
rect 3816 2799 3834 2826
rect 3942 2799 3960 2898
rect 3672 2754 3690 2781
rect 3762 2754 3780 2781
rect 3888 2754 3906 2781
rect 4131 2754 4149 2979
rect 4905 2880 4923 3276
rect 4689 2862 4923 2880
rect 4689 2835 4716 2862
rect 3654 2736 4149 2754
rect 4239 2817 4716 2835
rect 4239 2763 4257 2817
rect 4392 2763 4410 2817
rect 4689 2808 4716 2817
rect 4131 2583 4149 2736
rect 4293 2682 4311 2736
rect 4455 2682 4473 2745
rect 4761 2727 4788 2772
rect 4617 2691 4707 2718
rect 4761 2700 4815 2727
rect 4617 2682 4635 2691
rect 4293 2664 4635 2682
rect 4761 2682 4788 2700
rect 4410 2637 4419 2655
rect 4455 2628 4473 2664
rect 4689 2619 4716 2646
rect 4239 2583 4257 2601
rect 4689 2601 4788 2619
rect 4689 2583 4725 2601
rect 4131 2565 4725 2583
rect 4131 2052 4149 2565
rect 4905 2448 4923 2862
rect 4905 2430 5409 2448
rect 4905 2349 4923 2430
rect 4689 2331 4923 2349
rect 4689 2304 4716 2331
rect 4239 2286 4716 2304
rect 4239 2232 4257 2286
rect 4392 2232 4410 2286
rect 4689 2277 4716 2286
rect 4293 2151 4311 2205
rect 4455 2151 4473 2214
rect 4761 2196 4788 2241
rect 4617 2160 4707 2187
rect 4761 2169 4815 2196
rect 4617 2151 4635 2160
rect 4293 2133 4635 2151
rect 4761 2151 4788 2169
rect 4410 2106 4419 2124
rect 4455 2097 4473 2133
rect 4689 2088 4716 2115
rect 4239 2052 4257 2070
rect 4689 2070 4788 2088
rect 4689 2052 4725 2070
rect 3636 2034 4725 2052
rect 2223 1836 3213 1854
rect 2223 1071 2241 1836
rect 3186 1737 3213 1836
rect 3015 1719 3213 1737
rect 3015 1692 3042 1719
rect 2565 1674 3042 1692
rect 2565 1620 2583 1674
rect 2718 1620 2736 1674
rect 3015 1665 3042 1674
rect 2619 1539 2637 1593
rect 2781 1539 2799 1602
rect 2943 1548 3033 1575
rect 2943 1539 2961 1548
rect 2565 1512 2583 1530
rect 2619 1521 2961 1539
rect 3087 1539 3114 1629
rect 2718 1494 2736 1512
rect 2781 1485 2799 1521
rect 3015 1476 3042 1503
rect 2565 1440 2583 1458
rect 3015 1458 3114 1476
rect 3015 1440 3051 1458
rect 2475 1422 3051 1440
rect 2214 1053 2322 1071
rect 2223 1008 2250 1053
rect 2295 927 2322 972
rect 2475 972 2493 1422
rect 3186 1269 3213 1719
rect 3015 1251 3213 1269
rect 3015 1224 3042 1251
rect 2565 1206 3042 1224
rect 2565 1152 2583 1206
rect 2718 1152 2736 1206
rect 3015 1197 3042 1206
rect 2619 1071 2637 1125
rect 2781 1071 2799 1134
rect 3087 1116 3114 1161
rect 2943 1080 3033 1107
rect 3087 1089 3123 1116
rect 2943 1071 2961 1080
rect 2619 1053 2961 1071
rect 3087 1071 3114 1089
rect 2727 1026 2754 1044
rect 2781 1017 2799 1053
rect 3015 1008 3042 1035
rect 2565 972 2583 990
rect 3015 990 3114 1008
rect 3015 972 3051 990
rect 2475 954 3051 972
rect 2295 900 2340 927
rect 2295 882 2322 900
rect 2223 819 2250 846
rect 2475 819 2493 954
rect 3186 828 3213 1251
rect 2097 801 2493 819
rect 3015 810 3213 828
rect 2097 495 2115 801
rect 3015 783 3042 810
rect 2457 765 3042 783
rect 2457 756 2475 765
rect 2223 738 2475 756
rect 2223 729 2259 738
rect 2232 684 2259 729
rect 2565 711 2583 765
rect 2718 711 2736 765
rect 3015 756 3042 765
rect 2304 603 2331 648
rect 2619 630 2637 684
rect 2781 630 2799 693
rect 2943 639 3033 666
rect 2943 630 2961 639
rect 2565 612 2592 630
rect 2619 612 2961 630
rect 3087 630 3114 720
rect 2304 576 2367 603
rect 2781 576 2799 612
rect 2304 558 2331 576
rect 3015 567 3042 594
rect 2565 531 2583 549
rect 3015 549 3114 567
rect 3015 531 3051 549
rect 2232 495 2259 522
rect 2565 513 3051 531
rect 2565 495 2583 513
rect 2097 477 2583 495
rect 2232 117 2250 477
rect 3186 414 3213 810
rect 3015 396 3213 414
rect 3015 369 3042 396
rect 2565 351 3042 369
rect 2565 297 2583 351
rect 2718 297 2736 351
rect 3015 342 3042 351
rect 2619 216 2637 270
rect 2781 216 2799 279
rect 3087 261 3114 306
rect 2943 225 3033 252
rect 3087 234 3096 261
rect 2943 216 2961 225
rect 2619 198 2961 216
rect 3087 216 3114 234
rect 2781 162 2799 198
rect 3015 153 3042 180
rect 2565 117 2583 135
rect 3015 135 3114 153
rect 3015 117 3051 135
rect 2232 99 3051 117
rect 2862 -414 2880 99
rect 2925 45 2934 99
rect 3636 45 3654 2034
rect 5391 1818 5409 2430
rect 2925 27 3654 45
rect 4059 1800 5409 1818
rect 4059 -63 4077 1800
rect 5391 1701 5409 1800
rect 5490 1728 5724 1746
rect 5490 1701 5517 1728
rect 5040 1683 5517 1701
rect 5040 1629 5058 1683
rect 5193 1629 5211 1683
rect 5490 1674 5517 1683
rect 5094 1548 5112 1602
rect 5256 1548 5274 1611
rect 5562 1593 5589 1638
rect 5418 1557 5508 1584
rect 5562 1566 5616 1593
rect 5418 1548 5436 1557
rect 5094 1530 5436 1548
rect 5562 1548 5589 1566
rect 5202 1503 5220 1521
rect 5256 1494 5274 1530
rect 5490 1485 5517 1512
rect 5040 1449 5058 1467
rect 5490 1467 5589 1485
rect 5490 1449 5526 1467
rect 4932 1431 5526 1449
rect 4932 954 4950 1431
rect 5706 1251 5724 1728
rect 5490 1233 5724 1251
rect 5490 1206 5517 1233
rect 5040 1188 5517 1206
rect 5040 1134 5058 1188
rect 5193 1134 5211 1188
rect 5490 1179 5517 1188
rect 5094 1053 5112 1107
rect 5256 1053 5274 1116
rect 5562 1098 5589 1143
rect 5418 1062 5508 1089
rect 5562 1071 5616 1098
rect 5418 1053 5436 1062
rect 5094 1035 5436 1053
rect 5562 1053 5589 1071
rect 5193 1008 5220 1026
rect 5256 999 5274 1035
rect 5490 990 5517 1017
rect 5040 954 5058 972
rect 5490 972 5589 990
rect 5490 954 5526 972
rect 4932 936 5526 954
rect 4932 540 4950 936
rect 5706 837 5724 1233
rect 5490 819 5724 837
rect 5490 792 5517 819
rect 5040 774 5517 792
rect 5040 720 5058 774
rect 5193 720 5211 774
rect 5490 765 5517 774
rect 5094 639 5112 693
rect 5256 639 5274 702
rect 5562 684 5589 729
rect 5418 648 5508 675
rect 5562 657 5616 684
rect 5418 639 5436 648
rect 5094 621 5436 639
rect 5562 639 5589 657
rect 5202 594 5220 612
rect 5256 585 5274 621
rect 5490 576 5517 603
rect 5040 540 5058 558
rect 5490 558 5589 576
rect 5490 540 5526 558
rect 4932 522 5526 540
rect 4932 9 4950 522
rect 5706 306 5724 819
rect 5490 288 5724 306
rect 5490 261 5517 288
rect 5040 243 5517 261
rect 5040 189 5058 243
rect 5193 189 5211 243
rect 5490 234 5517 243
rect 5094 108 5112 162
rect 5256 108 5274 171
rect 5562 153 5589 198
rect 5418 117 5508 144
rect 5562 126 5616 153
rect 5418 108 5436 117
rect 5094 90 5436 108
rect 5562 108 5589 126
rect 5211 63 5220 81
rect 5256 54 5274 90
rect 5490 45 5517 72
rect 5706 54 5724 288
rect 6570 54 6588 63
rect 5040 9 5058 27
rect 5490 27 5589 45
rect 5706 36 6588 54
rect 5490 9 5526 27
rect 4932 -9 5526 9
rect 3879 -81 4113 -63
rect 3879 -108 3906 -81
rect 3429 -126 3906 -108
rect 3429 -180 3447 -126
rect 3582 -180 3600 -126
rect 3879 -135 3906 -126
rect 3483 -261 3501 -207
rect 3645 -261 3663 -198
rect 3807 -252 3897 -225
rect 3807 -261 3825 -252
rect 3483 -279 3825 -261
rect 3951 -261 3978 -171
rect 3582 -306 3609 -288
rect 3645 -315 3663 -279
rect 3879 -324 3906 -297
rect 3429 -360 3447 -342
rect 3879 -342 3978 -324
rect 3879 -360 3915 -342
rect 3321 -378 3915 -360
rect 3321 -414 3339 -378
rect 2862 -432 3339 -414
rect 3321 -855 3339 -432
rect 4095 -558 4113 -81
rect 5265 -315 5283 -9
rect 6570 -63 6588 36
rect 6669 -36 6903 -18
rect 6669 -63 6696 -36
rect 6219 -81 6696 -63
rect 6219 -135 6237 -81
rect 6372 -135 6390 -81
rect 6669 -90 6696 -81
rect 6273 -216 6291 -162
rect 6435 -216 6453 -153
rect 6741 -171 6768 -126
rect 6597 -207 6687 -180
rect 6741 -198 6795 -171
rect 6597 -216 6615 -207
rect 6273 -234 6615 -216
rect 6741 -216 6768 -198
rect 6381 -261 6399 -243
rect 6435 -270 6453 -234
rect 6669 -279 6696 -252
rect 6219 -315 6237 -297
rect 6669 -297 6768 -279
rect 6669 -315 6705 -297
rect 5265 -333 6705 -315
rect 3879 -576 4113 -558
rect 4401 -567 5211 -549
rect 3879 -603 3906 -576
rect 3429 -621 3906 -603
rect 3429 -675 3447 -621
rect 3582 -675 3600 -621
rect 3879 -630 3906 -621
rect 3483 -756 3501 -702
rect 3645 -756 3663 -693
rect 3807 -747 3897 -720
rect 3807 -756 3825 -747
rect 3483 -774 3825 -756
rect 3951 -756 3978 -666
rect 3591 -801 3600 -783
rect 3645 -810 3663 -774
rect 3879 -819 3906 -792
rect 3429 -855 3447 -837
rect 3879 -837 3978 -819
rect 3879 -855 3915 -837
rect 3321 -873 3915 -855
rect 3321 -1269 3339 -873
rect 4095 -972 4113 -576
rect 4491 -954 5022 -936
rect 3879 -990 4113 -972
rect 3879 -1017 3906 -990
rect 3429 -1035 3906 -1017
rect 3429 -1089 3447 -1035
rect 3582 -1089 3600 -1035
rect 3879 -1044 3906 -1035
rect 3483 -1170 3501 -1116
rect 3645 -1170 3663 -1107
rect 3951 -1125 3978 -1080
rect 3807 -1161 3897 -1134
rect 3951 -1152 3969 -1125
rect 3807 -1170 3825 -1161
rect 3483 -1188 3825 -1170
rect 3951 -1170 3978 -1152
rect 3645 -1224 3663 -1188
rect 3879 -1233 3906 -1206
rect 3429 -1269 3447 -1251
rect 3879 -1251 3978 -1233
rect 3879 -1269 3915 -1251
rect 3321 -1287 3915 -1269
rect 3321 -1773 3339 -1287
rect 4095 -1503 4113 -990
rect 4257 -1431 5148 -1413
rect 3879 -1521 4014 -1503
rect 3879 -1548 3906 -1521
rect 4032 -1521 4113 -1503
rect 3429 -1566 3906 -1548
rect 3429 -1620 3447 -1566
rect 3582 -1620 3600 -1566
rect 3879 -1575 3906 -1566
rect 3483 -1701 3501 -1647
rect 3645 -1701 3663 -1638
rect 3951 -1656 3978 -1611
rect 3807 -1692 3897 -1665
rect 3951 -1683 3969 -1656
rect 3807 -1701 3825 -1692
rect 3483 -1719 3825 -1701
rect 3951 -1701 3978 -1683
rect 3645 -1755 3663 -1719
rect 3276 -1791 3339 -1773
rect 3276 -2628 3294 -1791
rect 3321 -1800 3339 -1791
rect 3879 -1764 3906 -1737
rect 3429 -1800 3447 -1782
rect 3879 -1782 3978 -1764
rect 3879 -1800 3915 -1782
rect 3321 -1818 3915 -1800
rect 3726 -1881 3744 -1818
rect 5265 -1881 5283 -333
rect 5967 -378 6021 -360
rect 6111 -810 6129 -333
rect 6885 -513 6903 -36
rect 6669 -531 6903 -513
rect 6669 -558 6696 -531
rect 6219 -576 6696 -558
rect 6219 -630 6237 -576
rect 6372 -630 6390 -576
rect 6669 -585 6696 -576
rect 6273 -711 6291 -657
rect 6435 -711 6453 -648
rect 6741 -666 6768 -621
rect 6597 -702 6687 -675
rect 6741 -693 6795 -666
rect 6597 -711 6615 -702
rect 6273 -729 6615 -711
rect 6741 -711 6768 -693
rect 6372 -756 6399 -738
rect 6435 -765 6453 -729
rect 6669 -774 6696 -747
rect 6219 -810 6237 -792
rect 6669 -792 6768 -774
rect 6669 -810 6705 -792
rect 6111 -828 6705 -810
rect 5913 -927 6021 -909
rect 5913 -936 5931 -927
rect 6111 -1224 6129 -828
rect 6885 -927 6903 -531
rect 6669 -945 6903 -927
rect 6669 -972 6696 -945
rect 6219 -990 6696 -972
rect 6219 -1044 6237 -990
rect 6372 -1044 6390 -990
rect 6669 -999 6696 -990
rect 6273 -1125 6291 -1071
rect 6435 -1125 6453 -1062
rect 6741 -1080 6768 -1035
rect 6597 -1116 6687 -1089
rect 6741 -1107 6795 -1080
rect 6597 -1125 6615 -1116
rect 6273 -1143 6615 -1125
rect 6741 -1125 6768 -1107
rect 6381 -1170 6399 -1152
rect 6435 -1179 6453 -1143
rect 6669 -1188 6696 -1161
rect 6219 -1224 6237 -1206
rect 6669 -1206 6768 -1188
rect 6669 -1224 6705 -1206
rect 6111 -1242 6705 -1224
rect 6111 -1755 6129 -1242
rect 6885 -1458 6903 -945
rect 6669 -1476 6903 -1458
rect 6669 -1503 6696 -1476
rect 6219 -1521 6696 -1503
rect 6219 -1575 6237 -1521
rect 6372 -1575 6390 -1521
rect 6669 -1530 6696 -1521
rect 6273 -1656 6291 -1602
rect 6435 -1656 6453 -1593
rect 6741 -1611 6768 -1566
rect 6597 -1647 6687 -1620
rect 6741 -1638 6795 -1611
rect 6597 -1656 6615 -1647
rect 6273 -1674 6615 -1656
rect 6741 -1656 6768 -1638
rect 6390 -1701 6399 -1683
rect 6435 -1710 6453 -1674
rect 6669 -1719 6696 -1692
rect 6219 -1755 6237 -1737
rect 6669 -1737 6768 -1719
rect 6669 -1755 6705 -1737
rect 6111 -1773 6705 -1755
rect 3726 -1899 5283 -1881
rect 3519 -2241 3564 -2223
rect 4014 -2331 4032 -2169
rect 5544 -2232 5643 -2223
rect 5544 -2259 5571 -2232
rect 4932 -2277 5571 -2259
rect 4932 -2331 4950 -2277
rect 3834 -2349 4950 -2331
rect 5094 -2331 5112 -2277
rect 5247 -2331 5265 -2277
rect 5544 -2286 5571 -2277
rect 3834 -2376 3861 -2349
rect 3384 -2394 3861 -2376
rect 3384 -2448 3402 -2394
rect 3537 -2448 3555 -2394
rect 3834 -2403 3861 -2394
rect 3438 -2529 3456 -2475
rect 3600 -2529 3618 -2466
rect 3762 -2520 3852 -2493
rect 3906 -2502 3933 -2439
rect 3906 -2511 3960 -2502
rect 3762 -2529 3780 -2520
rect 3438 -2547 3780 -2529
rect 3906 -2529 3933 -2511
rect 3555 -2574 3573 -2556
rect 3600 -2583 3618 -2547
rect 3834 -2592 3861 -2565
rect 3384 -2628 3402 -2610
rect 3834 -2610 3933 -2592
rect 3834 -2628 3870 -2610
rect 3276 -2646 3870 -2628
rect 3276 -3123 3294 -2646
rect 3519 -2709 3528 -2691
rect 4050 -2826 4068 -2349
rect 4365 -2502 4851 -2484
rect 3834 -2844 4068 -2826
rect 3834 -2871 3861 -2844
rect 3384 -2889 3861 -2871
rect 3384 -2943 3402 -2889
rect 3537 -2943 3555 -2889
rect 3834 -2898 3861 -2889
rect 3438 -3024 3456 -2970
rect 3600 -3024 3618 -2961
rect 3906 -2979 3933 -2934
rect 3762 -3015 3852 -2988
rect 3906 -3006 3924 -2979
rect 3762 -3024 3780 -3015
rect 3438 -3042 3780 -3024
rect 3906 -3024 3933 -3006
rect 3546 -3069 3555 -3051
rect 3600 -3078 3618 -3042
rect 3834 -3087 3861 -3060
rect 3384 -3123 3402 -3105
rect 3834 -3105 3933 -3087
rect 3834 -3123 3870 -3105
rect 3276 -3141 3870 -3123
rect 3276 -3537 3294 -3141
rect 4050 -3240 4068 -2844
rect 3834 -3258 4068 -3240
rect 3834 -3285 3861 -3258
rect 3384 -3303 3861 -3285
rect 3384 -3357 3402 -3303
rect 3537 -3357 3555 -3303
rect 3834 -3312 3861 -3303
rect 3438 -3438 3456 -3384
rect 3600 -3438 3618 -3375
rect 3762 -3429 3852 -3402
rect 3762 -3438 3780 -3429
rect 3438 -3456 3780 -3438
rect 3906 -3438 3933 -3348
rect 3546 -3483 3564 -3465
rect 3600 -3492 3618 -3456
rect 3834 -3501 3861 -3474
rect 3384 -3537 3402 -3519
rect 3834 -3519 3933 -3501
rect 3834 -3537 3870 -3519
rect 3276 -3555 3870 -3537
rect 3276 -4068 3294 -3555
rect 4050 -3771 4068 -3258
rect 4932 -2736 4950 -2349
rect 5148 -2412 5166 -2358
rect 5310 -2412 5328 -2349
rect 5616 -2367 5643 -2322
rect 5472 -2403 5562 -2376
rect 5616 -2394 5670 -2367
rect 5472 -2412 5490 -2403
rect 5148 -2430 5490 -2412
rect 5616 -2412 5643 -2394
rect 5310 -2466 5328 -2430
rect 5544 -2475 5571 -2448
rect 5094 -2511 5112 -2493
rect 5544 -2493 5760 -2475
rect 5544 -2511 5580 -2493
rect 5094 -2529 5580 -2511
rect 5544 -2709 5643 -2700
rect 5544 -2736 5571 -2709
rect 4932 -2754 5571 -2736
rect 4932 -3132 4950 -2754
rect 5094 -2808 5112 -2754
rect 5247 -2808 5265 -2754
rect 5544 -2763 5571 -2754
rect 5148 -2889 5166 -2835
rect 5310 -2889 5328 -2826
rect 5616 -2844 5643 -2799
rect 5472 -2880 5562 -2853
rect 5616 -2871 5670 -2844
rect 5472 -2889 5490 -2880
rect 5148 -2907 5490 -2889
rect 5616 -2889 5643 -2871
rect 5310 -2943 5328 -2907
rect 5544 -2952 5571 -2925
rect 5742 -2952 5760 -2493
rect 5094 -2988 5112 -2970
rect 5544 -2970 5760 -2952
rect 5544 -2988 5580 -2970
rect 5094 -3006 5580 -2988
rect 5544 -3105 5643 -3096
rect 5544 -3132 5571 -3105
rect 4932 -3150 5571 -3132
rect 4932 -3600 4950 -3150
rect 5094 -3204 5112 -3150
rect 5247 -3204 5265 -3150
rect 5544 -3159 5571 -3150
rect 5148 -3285 5166 -3231
rect 5310 -3285 5328 -3222
rect 5616 -3240 5643 -3195
rect 5472 -3276 5562 -3249
rect 5616 -3267 5670 -3240
rect 5472 -3285 5490 -3276
rect 5148 -3303 5490 -3285
rect 5616 -3285 5643 -3267
rect 5256 -3330 5283 -3312
rect 5310 -3339 5328 -3303
rect 5544 -3348 5571 -3321
rect 5742 -3348 5760 -2970
rect 5094 -3384 5112 -3366
rect 5544 -3366 5760 -3348
rect 5544 -3384 5580 -3366
rect 5094 -3402 5580 -3384
rect 5544 -3573 5643 -3564
rect 5544 -3600 5571 -3573
rect 4932 -3618 5571 -3600
rect 5094 -3672 5112 -3618
rect 5247 -3672 5265 -3618
rect 5544 -3627 5571 -3618
rect 5148 -3753 5166 -3699
rect 5310 -3753 5328 -3690
rect 5616 -3708 5643 -3663
rect 5472 -3744 5562 -3717
rect 5616 -3735 5670 -3708
rect 5472 -3753 5490 -3744
rect 3834 -3789 4068 -3771
rect 4248 -3780 5067 -3762
rect 5148 -3771 5490 -3753
rect 5616 -3753 5643 -3735
rect 3834 -3816 3861 -3789
rect 3384 -3834 3861 -3816
rect 3384 -3888 3402 -3834
rect 3537 -3888 3555 -3834
rect 3834 -3843 3861 -3834
rect 3438 -3969 3456 -3915
rect 3600 -3969 3618 -3906
rect 3906 -3924 3933 -3879
rect 4248 -3924 4266 -3780
rect 5256 -3798 5283 -3780
rect 5310 -3807 5328 -3771
rect 5544 -3816 5571 -3789
rect 5742 -3816 5760 -3366
rect 5094 -3852 5112 -3834
rect 5544 -3834 5760 -3816
rect 5544 -3852 5580 -3834
rect 3762 -3960 3852 -3933
rect 3906 -3951 4266 -3924
rect 4932 -3870 5580 -3852
rect 3762 -3969 3780 -3960
rect 3438 -3987 3780 -3969
rect 3906 -3969 3933 -3951
rect 3555 -4014 3564 -3996
rect 3600 -4023 3618 -3987
rect 3834 -4032 3861 -4005
rect 3384 -4068 3402 -4050
rect 3834 -4050 3933 -4032
rect 3834 -4068 3870 -4050
rect 3276 -4086 3870 -4068
rect 3681 -4149 3699 -4086
rect 4932 -4149 4950 -3870
rect 3681 -4167 4950 -4149
<< m2contact >>
rect 4374 5490 4410 5508
rect 4356 4545 4410 4563
rect -279 4338 -216 4356
rect -45 4338 36 4356
rect 4374 3051 4410 3069
rect 4356 2106 4410 2124
rect 2520 1512 2565 1530
rect 2340 900 2367 927
rect 2520 612 2565 630
rect 5157 1008 5193 1026
rect 5184 63 5211 81
rect 3978 -738 4005 -711
rect 3546 -801 3591 -783
rect 4194 -1431 4257 -1413
rect 5148 -1431 5166 -1413
rect 3969 -1683 4005 -1656
rect 3555 -1746 3591 -1728
rect 6336 -756 6372 -738
rect 6021 -927 6057 -909
rect 6363 -1701 6390 -1683
rect 4671 -1935 4689 -1908
rect 3456 -2709 3519 -2691
rect 3501 -3069 3546 -3051
rect 5220 -3798 5256 -3780
rect 3519 -4014 3555 -3996
<< metal2 >>
rect -126 5823 4374 5841
rect -621 4338 -279 4356
rect -621 -4311 -603 4338
rect -126 -2691 -108 5823
rect 4356 5490 4374 5823
rect 4356 4356 4374 4545
rect 36 4338 4374 4356
rect 4356 3384 5337 3402
rect 4356 3051 4374 3384
rect 4356 1908 4374 2106
rect 738 1890 3645 1908
rect 3654 1890 4374 1908
rect 738 -2043 756 1890
rect 2385 1512 2520 1530
rect 2385 927 2403 1512
rect 5319 1350 5337 3384
rect 5157 1332 5337 1350
rect 5157 1026 5175 1332
rect 2367 900 2403 927
rect 2385 882 2403 900
rect 2385 864 2457 882
rect 2439 630 2457 864
rect 5157 855 5175 1008
rect 4671 837 5175 855
rect 2439 612 2520 630
rect 4671 -423 4689 837
rect 3546 -441 4689 -423
rect 5148 63 5184 81
rect 5211 63 5238 81
rect 3546 -783 3564 -441
rect 4005 -738 4689 -711
rect 3555 -1431 4194 -1413
rect 3555 -1728 3573 -1431
rect 4005 -1683 4131 -1656
rect 3555 -2043 3573 -1746
rect 738 -2061 3573 -2043
rect 4113 -2043 4131 -1683
rect 4671 -1908 4689 -738
rect 5148 -1413 5166 63
rect 6498 -414 6516 63
rect 6336 -432 6516 -414
rect 6336 -738 6354 -432
rect 6336 -909 6354 -756
rect 6057 -927 6354 -909
rect 6327 -1701 6363 -1683
rect 6390 -1701 6417 -1683
rect 4113 -2061 4752 -2043
rect -126 -2709 3456 -2691
rect 3501 -3051 3519 -2709
rect 4734 -3537 4752 -2061
rect 4734 -3555 5220 -3537
rect 5202 -3798 5220 -3555
rect 3510 -4014 3519 -3996
rect 3555 -4014 3582 -3996
rect 3510 -4311 3528 -4014
rect 6327 -4311 6345 -1701
rect -621 -4329 6345 -4311
<< m123contact >>
rect 4374 5985 4410 6003
rect -333 4878 -315 4896
rect 4374 5076 4410 5094
rect 378 4878 432 4896
rect 4131 4464 4149 4536
rect 4374 3546 4419 3564
rect 4131 3402 4149 3492
rect 4374 2637 4410 2655
rect 2682 1494 2718 1512
rect 5157 1503 5202 1521
rect 2673 1026 2727 1044
rect 2367 576 2421 603
rect 3546 -306 3582 -288
rect 5157 594 5202 612
rect 3969 -1152 4005 -1125
rect 3555 -1215 3591 -1197
rect 6336 -261 6381 -243
rect 6021 -378 6057 -360
rect 6336 -1170 6381 -1152
rect 3501 -2241 3519 -2223
rect 3501 -2574 3555 -2556
rect 3510 -3483 3546 -3465
rect 5229 -3330 5256 -3312
<< metal3 >>
rect 54 6291 4365 6318
rect -333 -3654 -315 4878
rect 54 -2178 72 6291
rect 4356 6003 4365 6291
rect 4356 5985 4374 6003
rect 4365 5076 4374 5094
rect 4365 4896 4383 5076
rect 432 4878 4383 4896
rect 4131 3492 4149 4464
rect 4356 3906 5175 3924
rect 4356 3546 4374 3906
rect 4365 2637 4374 2655
rect 4365 2457 4383 2637
rect 1224 2439 4383 2457
rect 1224 -1386 1242 2439
rect 5157 1521 5175 3906
rect 2682 1332 2700 1494
rect 5157 1404 5175 1503
rect 2403 1314 2700 1332
rect 4599 1386 5175 1404
rect 2403 945 2421 1314
rect 2673 945 2691 1026
rect 2403 927 2691 945
rect 2403 603 2421 927
rect 4599 81 4617 1386
rect 5157 441 5175 594
rect 3546 63 4617 81
rect 4752 423 5175 441
rect 3546 -288 3564 63
rect 4752 -891 4770 423
rect 6336 -243 6354 63
rect 6336 -360 6354 -261
rect 6057 -378 6354 -360
rect 3555 -909 4770 -891
rect 3555 -1197 3573 -909
rect 4005 -1152 4770 -1125
rect 3555 -1386 3573 -1215
rect 1224 -1404 3573 -1386
rect 4752 -1980 4770 -1152
rect 6336 -1323 6354 -1170
rect 4635 -1998 4770 -1980
rect 5940 -1341 6354 -1323
rect 54 -2205 3519 -2178
rect 3501 -2223 3519 -2205
rect 3501 -2556 3519 -2241
rect 4635 -3078 4653 -1998
rect 4635 -3096 5220 -3078
rect 5202 -3312 5220 -3096
rect 5202 -3330 5229 -3312
rect 3546 -3483 3564 -3465
rect 3510 -3636 3528 -3483
rect 3510 -3654 3519 -3636
rect -333 -3672 3519 -3654
rect 3024 -4464 3042 -3672
rect 5940 -4464 5958 -1341
rect 3024 -4482 5958 -4464
<< labels >>
rlabel polysilicon 2232 900 2232 900 1 s0
rlabel polysilicon 2223 576 2223 576 1 s1
rlabel m2contact 2358 909 2358 909 1 s0_not
rlabel metal1 2358 594 2358 594 1 s1_not
rlabel polysilicon 3276 1566 3276 1566 1 D0
rlabel polysilicon 3258 1107 3258 1107 1 D1
rlabel polysilicon 3249 666 3249 666 1 D2
rlabel polysilicon 3195 252 3195 252 1 D3
rlabel metal3 3555 -54 3555 -54 1 a3
rlabel metal2 3555 -531 3555 -531 1 a2
rlabel metal3 3564 -1341 3564 -1341 1 a1
rlabel metal2 3564 -1899 3564 -1899 1 a0
rlabel metal2 3519 -4149 3519 -4149 1 b0
rlabel metal3 3519 -3618 3519 -3618 1 b1
rlabel metal2 3510 -2817 3510 -2817 1 b2
rlabel metal3 3510 -2304 3510 -2304 1 b3
rlabel metal1 3933 -3933 3933 -3933 1 and_b0
rlabel polycontact 3951 -3402 3951 -3402 1 and_b1
rlabel polycontact 3942 -2988 3942 -2988 1 and_b2
rlabel metal1 3942 -2502 3942 -2502 1 and_b3
rlabel metal1 3978 -234 3978 -234 1 and_a3
rlabel metal1 3969 -1674 3969 -1674 1 and_a0
rlabel m123contact 3978 -1143 3978 -1143 1 and_a1
rlabel metal1 3978 -729 3978 -729 1 and_a2
rlabel metal1 5643 -3717 5643 -3717 1 and_oper_out0
rlabel metal1 5643 -3249 5643 -3249 1 and_oper_out1
rlabel metal1 5652 -2862 5652 -2862 1 and_oper_out2
rlabel metal1 5652 -2385 5652 -2385 1 and_oper_out3
rlabel metal1 5598 1080 5598 1080 1 comp_a2
rlabel metal1 5598 1584 5598 1584 1 comp_a3
rlabel metal1 5589 675 5589 675 1 comp_a1
rlabel metal1 5598 135 5598 135 1 comp_a0
rlabel metal1 6768 -189 6768 -189 1 comp_b3
rlabel metal1 6759 -684 6759 -684 1 comp_b2
rlabel metal1 6768 -1098 6768 -1098 1 comp_b1
rlabel metal1 6777 -1629 6777 -1629 1 comp_b0
rlabel metal1 4797 2178 4797 2178 1 adsub_a0
rlabel metal1 4797 2709 4797 2709 1 adsub_a1
rlabel metal1 4788 3123 4788 3123 1 adsub_a2
rlabel metal1 4788 3618 4788 3618 1 adsub_a3
rlabel metal1 4797 6057 4797 6057 1 adsub_b3
rlabel metal1 4806 5571 4806 5571 1 adsub_b2
rlabel metal1 4797 5148 4797 5148 1 adsub_b1
rlabel metal1 4797 4626 4797 4626 1 adsub_b0
<< end >>
