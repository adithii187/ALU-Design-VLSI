magic
tech scmos
timestamp 1700396393
<< nwell >>
rect 279 1080 1260 1098
rect 1035 981 1224 1008
rect 1233 981 1260 1080
rect 1035 963 1260 981
rect 1035 954 1224 963
rect 567 801 891 891
rect 1035 846 1188 954
rect 1035 837 1098 846
rect 1116 837 1188 846
rect 1035 513 1224 540
rect 1233 513 1260 963
rect 1035 495 1260 513
rect 1035 486 1224 495
rect 234 315 423 342
rect 567 333 891 423
rect 1035 378 1188 486
rect 1035 369 1098 378
rect 1116 369 1188 378
rect 234 297 261 315
rect 369 297 423 315
rect 243 189 396 297
rect 243 180 306 189
rect 324 180 396 189
rect 1035 72 1224 99
rect 1233 72 1260 495
rect 1035 54 1260 72
rect 1035 45 1224 54
rect 243 0 432 18
rect 504 0 522 27
rect 243 -18 522 0
rect 243 -27 432 -18
rect 252 -135 405 -27
rect 567 -108 891 -18
rect 1035 -63 1188 45
rect 1035 -72 1098 -63
rect 1116 -72 1188 -63
rect 252 -144 315 -135
rect 333 -144 405 -135
rect 1035 -342 1224 -315
rect 1233 -342 1260 54
rect 1035 -360 1260 -342
rect 1035 -369 1224 -360
rect 567 -522 891 -432
rect 1035 -477 1188 -369
rect 1035 -486 1098 -477
rect 1116 -486 1188 -477
<< ntransistor >>
rect 1098 756 1116 783
rect 639 702 657 729
rect 801 702 819 729
rect 1098 288 1116 315
rect 639 234 657 261
rect 801 234 819 261
rect 306 99 324 126
rect 1098 -153 1116 -126
rect 315 -225 333 -198
rect 639 -207 657 -180
rect 774 -207 792 -180
rect 801 -207 819 -180
rect 1098 -567 1116 -540
rect 639 -621 657 -594
rect 756 -621 774 -594
rect 801 -621 819 -594
<< ptransistor >>
rect 639 828 657 873
rect 801 828 819 873
rect 1098 855 1116 909
rect 639 360 657 405
rect 801 360 819 405
rect 1098 387 1116 441
rect 306 198 324 252
rect 315 -126 333 -72
rect 639 -81 657 -36
rect 801 -81 819 -36
rect 1098 -54 1116 0
rect 639 -495 657 -450
rect 801 -495 819 -450
rect 1098 -468 1116 -414
<< ndiffusion >>
rect 1053 774 1098 783
rect 1053 756 1062 774
rect 1089 756 1098 774
rect 1116 756 1134 783
rect 1161 756 1170 783
rect 603 720 639 729
rect 603 702 612 720
rect 630 702 639 720
rect 657 702 801 729
rect 819 711 828 729
rect 846 711 855 729
rect 819 702 855 711
rect 1053 306 1098 315
rect 1053 288 1062 306
rect 1089 288 1098 306
rect 1116 288 1134 315
rect 1161 288 1170 315
rect 603 252 639 261
rect 603 234 612 252
rect 630 234 639 252
rect 657 234 801 261
rect 819 243 828 261
rect 846 243 855 261
rect 819 234 855 243
rect 261 117 306 126
rect 261 99 270 117
rect 297 99 306 117
rect 324 99 342 126
rect 369 99 378 126
rect 1053 -135 1098 -126
rect 1053 -153 1062 -135
rect 1089 -153 1098 -135
rect 1116 -153 1134 -126
rect 1161 -153 1170 -126
rect 603 -189 639 -180
rect 270 -207 315 -198
rect 270 -225 279 -207
rect 306 -225 315 -207
rect 333 -225 351 -198
rect 378 -225 387 -198
rect 603 -207 612 -189
rect 630 -207 639 -189
rect 657 -207 774 -180
rect 792 -207 801 -180
rect 819 -198 828 -180
rect 846 -198 855 -180
rect 819 -207 855 -198
rect 1053 -549 1098 -540
rect 1053 -567 1062 -549
rect 1089 -567 1098 -549
rect 1116 -567 1134 -540
rect 1161 -567 1170 -540
rect 603 -603 639 -594
rect 603 -621 612 -603
rect 630 -621 639 -603
rect 657 -621 756 -594
rect 774 -621 801 -594
rect 819 -612 828 -594
rect 846 -612 855 -594
rect 819 -621 855 -612
<< pdiffusion >>
rect 1053 882 1062 909
rect 1089 882 1098 909
rect 603 864 639 873
rect 603 846 612 864
rect 630 846 639 864
rect 603 828 639 846
rect 657 855 720 873
rect 657 837 666 855
rect 684 837 720 855
rect 657 828 720 837
rect 756 864 801 873
rect 756 846 765 864
rect 783 846 801 864
rect 756 828 801 846
rect 819 864 855 873
rect 819 846 828 864
rect 846 846 855 864
rect 1053 855 1098 882
rect 1116 900 1170 909
rect 1116 873 1134 900
rect 1161 873 1170 900
rect 1116 855 1170 873
rect 819 828 855 846
rect 1053 414 1062 441
rect 1089 414 1098 441
rect 603 396 639 405
rect 603 378 612 396
rect 630 378 639 396
rect 603 360 639 378
rect 657 387 720 405
rect 657 369 666 387
rect 684 369 720 387
rect 657 360 720 369
rect 756 396 801 405
rect 756 378 765 396
rect 783 378 801 396
rect 756 360 801 378
rect 819 396 855 405
rect 819 378 828 396
rect 846 378 855 396
rect 1053 387 1098 414
rect 1116 432 1170 441
rect 1116 405 1134 432
rect 1161 405 1170 432
rect 1116 387 1170 405
rect 819 360 855 378
rect 261 225 270 252
rect 297 225 306 252
rect 261 198 306 225
rect 324 243 378 252
rect 324 216 342 243
rect 369 216 378 243
rect 324 198 378 216
rect 1053 -27 1062 0
rect 1089 -27 1098 0
rect 603 -45 639 -36
rect 603 -63 612 -45
rect 630 -63 639 -45
rect 270 -99 279 -72
rect 306 -99 315 -72
rect 270 -126 315 -99
rect 333 -81 387 -72
rect 603 -81 639 -63
rect 657 -54 720 -36
rect 657 -72 666 -54
rect 684 -72 720 -54
rect 657 -81 720 -72
rect 756 -45 801 -36
rect 756 -63 765 -45
rect 783 -63 801 -45
rect 756 -81 801 -63
rect 819 -45 855 -36
rect 819 -63 828 -45
rect 846 -63 855 -45
rect 1053 -54 1098 -27
rect 1116 -9 1170 0
rect 1116 -36 1134 -9
rect 1161 -36 1170 -9
rect 1116 -54 1170 -36
rect 819 -81 855 -63
rect 333 -108 351 -81
rect 378 -108 387 -81
rect 333 -126 387 -108
rect 1053 -441 1062 -414
rect 1089 -441 1098 -414
rect 603 -459 639 -450
rect 603 -477 612 -459
rect 630 -477 639 -459
rect 603 -495 639 -477
rect 657 -468 720 -450
rect 657 -486 666 -468
rect 684 -486 720 -468
rect 657 -495 720 -486
rect 756 -459 801 -450
rect 756 -477 765 -459
rect 783 -477 801 -459
rect 756 -495 801 -477
rect 819 -459 855 -450
rect 819 -477 828 -459
rect 846 -477 855 -459
rect 1053 -468 1098 -441
rect 1116 -423 1170 -414
rect 1116 -450 1134 -423
rect 1161 -450 1170 -423
rect 1116 -468 1170 -450
rect 819 -495 855 -477
<< ndcontact >>
rect 1062 747 1089 774
rect 1134 756 1161 783
rect 612 702 630 720
rect 828 711 846 729
rect 1062 279 1089 306
rect 1134 288 1161 315
rect 612 234 630 252
rect 828 243 846 261
rect 270 90 297 117
rect 342 99 369 126
rect 1062 -162 1089 -135
rect 1134 -153 1161 -126
rect 279 -234 306 -207
rect 351 -225 378 -198
rect 612 -207 630 -189
rect 828 -198 846 -180
rect 1062 -576 1089 -549
rect 1134 -567 1161 -540
rect 612 -621 630 -603
rect 828 -612 846 -594
<< pdcontact >>
rect 1062 882 1089 909
rect 612 846 630 864
rect 666 837 684 855
rect 765 846 783 864
rect 828 846 846 864
rect 1134 873 1161 900
rect 1062 414 1089 441
rect 612 378 630 396
rect 666 369 684 387
rect 765 378 783 396
rect 828 378 846 396
rect 1134 405 1161 432
rect 270 225 297 252
rect 342 216 369 243
rect 1062 -27 1089 0
rect 612 -63 630 -45
rect 279 -99 306 -72
rect 666 -72 684 -54
rect 765 -63 783 -45
rect 828 -63 846 -45
rect 1134 -36 1161 -9
rect 351 -108 378 -81
rect 1062 -441 1089 -414
rect 612 -477 630 -459
rect 666 -486 684 -468
rect 765 -477 783 -459
rect 828 -477 846 -459
rect 1134 -450 1161 -423
<< polysilicon >>
rect 1098 909 1116 1026
rect 639 873 657 900
rect 801 873 819 900
rect 639 774 657 828
rect 801 756 819 828
rect 1098 819 1116 855
rect 1107 792 1116 819
rect 1098 783 1116 792
rect 639 729 657 756
rect 1098 738 1116 756
rect 801 729 819 738
rect 639 693 657 702
rect 801 693 819 702
rect 171 441 567 459
rect 1098 441 1116 558
rect 171 162 189 441
rect 549 297 567 441
rect 639 405 657 432
rect 801 405 819 432
rect 639 297 657 360
rect 549 279 657 297
rect 306 252 324 270
rect 639 261 657 279
rect 801 288 819 360
rect 1098 351 1116 387
rect 1107 324 1116 351
rect 1098 315 1116 324
rect 1098 270 1116 288
rect 801 261 819 270
rect 639 225 657 234
rect 801 225 819 234
rect 306 162 324 198
rect 54 135 324 162
rect 54 -702 72 135
rect 306 126 324 135
rect 306 81 324 99
rect 1098 0 1116 117
rect 639 -36 657 -9
rect 801 -36 819 -9
rect 315 -72 333 -54
rect 639 -126 657 -81
rect 315 -162 333 -126
rect 108 -189 333 -162
rect 639 -180 657 -144
rect 801 -153 819 -81
rect 1098 -90 1116 -54
rect 1107 -117 1116 -90
rect 1098 -126 1116 -117
rect 774 -171 819 -153
rect 1098 -171 1116 -153
rect 774 -180 792 -171
rect 801 -180 819 -171
rect 108 -306 126 -189
rect 315 -198 333 -189
rect 639 -216 657 -207
rect 315 -243 333 -225
rect 774 -306 792 -207
rect 801 -216 819 -207
rect 108 -324 792 -306
rect 495 -531 513 -324
rect 1098 -414 1116 -297
rect 639 -450 657 -423
rect 801 -450 819 -423
rect 639 -531 657 -495
rect 495 -549 657 -531
rect 639 -594 657 -549
rect 801 -567 819 -495
rect 1098 -504 1116 -468
rect 1107 -531 1116 -504
rect 1098 -540 1116 -531
rect 756 -585 819 -567
rect 1098 -585 1116 -567
rect 756 -594 774 -585
rect 801 -594 819 -585
rect 639 -630 657 -621
rect 756 -702 774 -621
rect 801 -630 819 -621
rect 54 -720 774 -702
<< polycontact >>
rect 630 756 657 774
rect 1080 792 1107 819
rect 783 738 819 756
rect 1080 324 1107 351
rect 801 270 819 288
rect 639 -144 657 -126
rect 1080 -117 1107 -90
rect 1080 -531 1107 -504
<< metal1 >>
rect 270 1080 1260 1098
rect 270 315 288 1080
rect 1233 981 1260 1080
rect 1062 963 1260 981
rect 1062 936 1089 963
rect 612 918 1089 936
rect 612 864 630 918
rect 765 864 783 918
rect 1062 909 1089 918
rect 666 783 684 837
rect 828 783 846 846
rect 1134 828 1161 873
rect 990 792 1080 819
rect 1134 801 1188 828
rect 990 783 1008 792
rect 612 756 630 774
rect 666 765 1008 783
rect 1134 783 1161 801
rect 765 738 783 756
rect 828 729 846 765
rect 1062 720 1089 747
rect 612 684 630 702
rect 1062 702 1161 720
rect 1062 684 1098 702
rect 522 666 1098 684
rect 261 297 369 315
rect 270 252 297 297
rect 342 171 369 216
rect 522 216 540 666
rect 1233 513 1260 963
rect 1062 495 1260 513
rect 1062 468 1089 495
rect 612 450 1089 468
rect 612 396 630 450
rect 765 396 783 450
rect 1062 441 1089 450
rect 666 315 684 369
rect 828 315 846 378
rect 1134 360 1161 405
rect 990 324 1080 351
rect 1134 333 1188 360
rect 990 315 1008 324
rect 666 297 1008 315
rect 1134 315 1161 333
rect 774 270 801 288
rect 828 261 846 297
rect 1062 252 1089 279
rect 612 216 630 234
rect 1062 234 1161 252
rect 1062 216 1098 234
rect 522 198 1098 216
rect 342 144 423 171
rect 342 126 369 144
rect 270 63 297 90
rect 522 63 540 198
rect 1233 72 1260 495
rect 144 45 540 63
rect 1062 54 1260 72
rect 144 -261 162 45
rect 1062 27 1089 54
rect 504 9 1089 27
rect 504 0 522 9
rect 270 -18 522 0
rect 270 -27 306 -18
rect 279 -72 306 -27
rect 612 -45 630 9
rect 765 -45 783 9
rect 1062 0 1089 9
rect 351 -153 378 -108
rect 666 -126 684 -72
rect 828 -126 846 -63
rect 1134 -81 1161 -36
rect 990 -117 1080 -90
rect 1134 -108 1188 -81
rect 990 -126 1008 -117
rect 603 -144 639 -126
rect 666 -144 1008 -126
rect 1134 -126 1161 -108
rect 351 -180 414 -153
rect 828 -180 846 -144
rect 351 -198 378 -180
rect 1062 -189 1089 -162
rect 612 -225 630 -207
rect 1062 -207 1161 -189
rect 1062 -225 1098 -207
rect 279 -261 306 -234
rect 612 -243 1098 -225
rect 612 -261 630 -243
rect 144 -279 630 -261
rect 279 -639 297 -279
rect 1233 -342 1260 54
rect 1062 -360 1260 -342
rect 1062 -387 1089 -360
rect 612 -405 1089 -387
rect 612 -459 630 -405
rect 765 -459 783 -405
rect 1062 -414 1089 -405
rect 666 -540 684 -486
rect 828 -540 846 -477
rect 1134 -495 1161 -450
rect 990 -531 1080 -504
rect 1134 -522 1188 -495
rect 990 -540 1008 -531
rect 666 -558 1008 -540
rect 1134 -540 1161 -522
rect 828 -594 846 -558
rect 1062 -603 1089 -576
rect 612 -639 630 -621
rect 1062 -621 1161 -603
rect 1062 -639 1098 -621
rect 279 -657 1098 -639
<< m2contact >>
rect 567 756 612 774
rect 423 144 450 171
rect 567 -144 603 -126
<< metal2 >>
rect 432 756 567 774
rect 432 171 450 756
rect 450 144 504 171
rect 486 -126 504 144
rect 486 -144 567 -126
<< m123contact >>
rect 729 738 765 756
rect 720 270 774 288
rect 414 -180 468 -153
<< metal3 >>
rect 729 576 747 738
rect 450 558 747 576
rect 450 189 468 558
rect 720 189 738 270
rect 450 171 738 189
rect 450 -153 468 171
<< labels >>
rlabel polysilicon 180 225 180 225 1 s0
rlabel polysilicon 234 -171 234 -171 1 s1
rlabel metal1 279 621 279 621 1 vdd
rlabel metal1 396 -648 396 -648 1 gnd
rlabel metal1 1179 -513 1179 -513 1 D3
rlabel metal1 1179 -99 1179 -99 1 D2
rlabel metal1 1161 342 1161 342 1 D1
rlabel metal1 1170 819 1170 819 1 D0
rlabel metal1 396 153 396 153 1 s0_not
rlabel metal1 405 -171 405 -171 1 s1_not
<< end >>
