magic
tech scmos
timestamp 1701322998
<< nwell >>
rect 477 -1728 585 -1053
rect 1287 -1728 1395 -1053
rect 2169 -1728 2277 -1053
rect 1827 -1917 2016 -1863
rect 801 -1980 990 -1926
rect 333 -2133 657 -2043
rect 801 -2088 954 -1980
rect 1359 -2070 1683 -1980
rect 1827 -2025 1980 -1917
rect 1827 -2034 1890 -2025
rect 1908 -2034 1980 -2025
rect 801 -2097 864 -2088
rect 882 -2097 954 -2088
rect 1017 -2484 1368 -2367
rect 477 -3825 585 -3150
rect 1287 -3825 1395 -3150
rect 2169 -3825 2277 -3150
rect 1827 -4014 2016 -3960
rect 801 -4077 990 -4023
rect 333 -4230 657 -4140
rect 801 -4185 954 -4077
rect 1359 -4167 1683 -4077
rect 1827 -4122 1980 -4014
rect 1827 -4131 1890 -4122
rect 1908 -4131 1980 -4122
rect 801 -4194 864 -4185
rect 882 -4194 954 -4185
rect 1017 -4581 1368 -4464
rect 477 -5940 585 -5265
rect 1287 -5940 1395 -5265
rect 2169 -5940 2277 -5265
rect 1827 -6129 2016 -6075
rect 801 -6192 990 -6138
rect 333 -6345 657 -6255
rect 801 -6300 954 -6192
rect 1359 -6282 1683 -6192
rect 1827 -6237 1980 -6129
rect 1827 -6246 1890 -6237
rect 1908 -6246 1980 -6237
rect 801 -6309 864 -6300
rect 882 -6309 954 -6300
rect 1017 -6696 1368 -6579
rect 477 -7875 585 -7200
rect 1287 -7875 1395 -7200
rect 2169 -7875 2277 -7200
rect 1827 -8064 2016 -8010
rect 801 -8127 990 -8073
rect 333 -8280 657 -8190
rect 801 -8235 954 -8127
rect 1359 -8217 1683 -8127
rect 1827 -8172 1980 -8064
rect 1827 -8181 1890 -8172
rect 1908 -8181 1980 -8172
rect 801 -8244 864 -8235
rect 882 -8244 954 -8235
rect 1017 -8631 1368 -8514
<< ntransistor >>
rect 252 -1134 306 -1116
rect 1062 -1134 1116 -1116
rect 252 -1305 306 -1287
rect 252 -1503 306 -1485
rect 252 -1665 306 -1647
rect 1944 -1134 1998 -1116
rect 1062 -1305 1116 -1287
rect 1062 -1503 1116 -1485
rect 1062 -1665 1116 -1647
rect 1944 -1305 1998 -1287
rect 1944 -1503 1998 -1485
rect 1944 -1665 1998 -1647
rect 864 -2178 882 -2151
rect 405 -2232 423 -2205
rect 567 -2232 585 -2205
rect 1431 -2169 1449 -2142
rect 1593 -2169 1611 -2142
rect 1890 -2115 1908 -2088
rect 1080 -2583 1098 -2556
rect 1170 -2583 1188 -2556
rect 1296 -2583 1314 -2556
rect 252 -3231 306 -3213
rect 1062 -3231 1116 -3213
rect 252 -3402 306 -3384
rect 252 -3600 306 -3582
rect 252 -3762 306 -3744
rect 1944 -3231 1998 -3213
rect 1062 -3402 1116 -3384
rect 1062 -3600 1116 -3582
rect 1062 -3762 1116 -3744
rect 1944 -3402 1998 -3384
rect 1944 -3600 1998 -3582
rect 1944 -3762 1998 -3744
rect 864 -4275 882 -4248
rect 405 -4329 423 -4302
rect 567 -4329 585 -4302
rect 1431 -4266 1449 -4239
rect 1593 -4266 1611 -4239
rect 1890 -4212 1908 -4185
rect 1080 -4680 1098 -4653
rect 1170 -4680 1188 -4653
rect 1296 -4680 1314 -4653
rect 252 -5346 306 -5328
rect 1062 -5346 1116 -5328
rect 252 -5517 306 -5499
rect 252 -5715 306 -5697
rect 252 -5877 306 -5859
rect 1944 -5346 1998 -5328
rect 1062 -5517 1116 -5499
rect 1062 -5715 1116 -5697
rect 1062 -5877 1116 -5859
rect 1944 -5517 1998 -5499
rect 1944 -5715 1998 -5697
rect 1944 -5877 1998 -5859
rect 864 -6390 882 -6363
rect 405 -6444 423 -6417
rect 567 -6444 585 -6417
rect 1431 -6381 1449 -6354
rect 1593 -6381 1611 -6354
rect 1890 -6327 1908 -6300
rect 1080 -6795 1098 -6768
rect 1170 -6795 1188 -6768
rect 1296 -6795 1314 -6768
rect 252 -7281 306 -7263
rect 1062 -7281 1116 -7263
rect 252 -7452 306 -7434
rect 252 -7650 306 -7632
rect 252 -7812 306 -7794
rect 1944 -7281 1998 -7263
rect 1062 -7452 1116 -7434
rect 1062 -7650 1116 -7632
rect 1062 -7812 1116 -7794
rect 1944 -7452 1998 -7434
rect 1944 -7650 1998 -7632
rect 1944 -7812 1998 -7794
rect 864 -8325 882 -8298
rect 405 -8379 423 -8352
rect 567 -8379 585 -8352
rect 1431 -8316 1449 -8289
rect 1593 -8316 1611 -8289
rect 1890 -8262 1908 -8235
rect 1080 -8730 1098 -8703
rect 1170 -8730 1188 -8703
rect 1296 -8730 1314 -8703
<< ptransistor >>
rect 504 -1134 567 -1116
rect 1314 -1134 1377 -1116
rect 504 -1305 567 -1287
rect 504 -1503 567 -1485
rect 504 -1665 567 -1647
rect 2196 -1134 2259 -1116
rect 1314 -1305 1377 -1287
rect 1314 -1503 1377 -1485
rect 1314 -1665 1377 -1647
rect 2196 -1305 2259 -1287
rect 2196 -1503 2259 -1485
rect 2196 -1665 2259 -1647
rect 405 -2106 423 -2061
rect 567 -2106 585 -2061
rect 864 -2079 882 -2025
rect 1431 -2043 1449 -1998
rect 1593 -2043 1611 -1998
rect 1890 -2016 1908 -1962
rect 1080 -2466 1098 -2421
rect 1170 -2466 1188 -2421
rect 1296 -2466 1314 -2421
rect 504 -3231 567 -3213
rect 1314 -3231 1377 -3213
rect 504 -3402 567 -3384
rect 504 -3600 567 -3582
rect 504 -3762 567 -3744
rect 2196 -3231 2259 -3213
rect 1314 -3402 1377 -3384
rect 1314 -3600 1377 -3582
rect 1314 -3762 1377 -3744
rect 2196 -3402 2259 -3384
rect 2196 -3600 2259 -3582
rect 2196 -3762 2259 -3744
rect 405 -4203 423 -4158
rect 567 -4203 585 -4158
rect 864 -4176 882 -4122
rect 1431 -4140 1449 -4095
rect 1593 -4140 1611 -4095
rect 1890 -4113 1908 -4059
rect 1080 -4563 1098 -4518
rect 1170 -4563 1188 -4518
rect 1296 -4563 1314 -4518
rect 504 -5346 567 -5328
rect 1314 -5346 1377 -5328
rect 504 -5517 567 -5499
rect 504 -5715 567 -5697
rect 504 -5877 567 -5859
rect 2196 -5346 2259 -5328
rect 1314 -5517 1377 -5499
rect 1314 -5715 1377 -5697
rect 1314 -5877 1377 -5859
rect 2196 -5517 2259 -5499
rect 2196 -5715 2259 -5697
rect 2196 -5877 2259 -5859
rect 405 -6318 423 -6273
rect 567 -6318 585 -6273
rect 864 -6291 882 -6237
rect 1431 -6255 1449 -6210
rect 1593 -6255 1611 -6210
rect 1890 -6228 1908 -6174
rect 1080 -6678 1098 -6633
rect 1170 -6678 1188 -6633
rect 1296 -6678 1314 -6633
rect 504 -7281 567 -7263
rect 1314 -7281 1377 -7263
rect 504 -7452 567 -7434
rect 504 -7650 567 -7632
rect 504 -7812 567 -7794
rect 2196 -7281 2259 -7263
rect 1314 -7452 1377 -7434
rect 1314 -7650 1377 -7632
rect 1314 -7812 1377 -7794
rect 2196 -7452 2259 -7434
rect 2196 -7650 2259 -7632
rect 2196 -7812 2259 -7794
rect 405 -8253 423 -8208
rect 567 -8253 585 -8208
rect 864 -8226 882 -8172
rect 1431 -8190 1449 -8145
rect 1593 -8190 1611 -8145
rect 1890 -8163 1908 -8109
rect 1080 -8613 1098 -8568
rect 1170 -8613 1188 -8568
rect 1296 -8613 1314 -8568
<< ndiffusion >>
rect 252 -1071 306 -1062
rect 252 -1107 261 -1071
rect 297 -1107 306 -1071
rect 252 -1116 306 -1107
rect 252 -1143 306 -1134
rect 252 -1179 261 -1143
rect 297 -1179 306 -1143
rect 252 -1188 306 -1179
rect 252 -1242 306 -1233
rect 252 -1278 261 -1242
rect 297 -1278 306 -1242
rect 252 -1287 306 -1278
rect 1062 -1071 1116 -1062
rect 1062 -1107 1071 -1071
rect 1107 -1107 1116 -1071
rect 1062 -1116 1116 -1107
rect 252 -1314 306 -1305
rect 252 -1350 261 -1314
rect 297 -1350 306 -1314
rect 252 -1359 306 -1350
rect 252 -1431 306 -1422
rect 252 -1467 261 -1431
rect 297 -1467 306 -1431
rect 252 -1485 306 -1467
rect 252 -1512 306 -1503
rect 252 -1548 261 -1512
rect 297 -1548 306 -1512
rect 252 -1557 306 -1548
rect 252 -1593 306 -1584
rect 252 -1629 261 -1593
rect 297 -1629 306 -1593
rect 252 -1647 306 -1629
rect 252 -1674 306 -1665
rect 252 -1710 261 -1674
rect 297 -1710 306 -1674
rect 252 -1719 306 -1710
rect 1062 -1143 1116 -1134
rect 1062 -1179 1071 -1143
rect 1107 -1179 1116 -1143
rect 1062 -1188 1116 -1179
rect 1062 -1242 1116 -1233
rect 1062 -1278 1071 -1242
rect 1107 -1278 1116 -1242
rect 1062 -1287 1116 -1278
rect 1944 -1071 1998 -1062
rect 1944 -1107 1953 -1071
rect 1989 -1107 1998 -1071
rect 1944 -1116 1998 -1107
rect 1062 -1314 1116 -1305
rect 1062 -1350 1071 -1314
rect 1107 -1350 1116 -1314
rect 1062 -1359 1116 -1350
rect 1062 -1431 1116 -1422
rect 1062 -1467 1071 -1431
rect 1107 -1467 1116 -1431
rect 1062 -1485 1116 -1467
rect 1062 -1512 1116 -1503
rect 1062 -1548 1071 -1512
rect 1107 -1548 1116 -1512
rect 1062 -1557 1116 -1548
rect 1062 -1593 1116 -1584
rect 1062 -1629 1071 -1593
rect 1107 -1629 1116 -1593
rect 1062 -1647 1116 -1629
rect 1062 -1674 1116 -1665
rect 1062 -1710 1071 -1674
rect 1107 -1710 1116 -1674
rect 1062 -1719 1116 -1710
rect 1944 -1143 1998 -1134
rect 1944 -1179 1953 -1143
rect 1989 -1179 1998 -1143
rect 1944 -1188 1998 -1179
rect 1944 -1242 1998 -1233
rect 1944 -1278 1953 -1242
rect 1989 -1278 1998 -1242
rect 1944 -1287 1998 -1278
rect 1944 -1314 1998 -1305
rect 1944 -1350 1953 -1314
rect 1989 -1350 1998 -1314
rect 1944 -1359 1998 -1350
rect 1944 -1431 1998 -1422
rect 1944 -1467 1953 -1431
rect 1989 -1467 1998 -1431
rect 1944 -1485 1998 -1467
rect 1944 -1512 1998 -1503
rect 1944 -1548 1953 -1512
rect 1989 -1548 1998 -1512
rect 1944 -1557 1998 -1548
rect 1944 -1593 1998 -1584
rect 1944 -1629 1953 -1593
rect 1989 -1629 1998 -1593
rect 1944 -1647 1998 -1629
rect 1944 -1674 1998 -1665
rect 1944 -1710 1953 -1674
rect 1989 -1710 1998 -1674
rect 1944 -1719 1998 -1710
rect 819 -2160 864 -2151
rect 819 -2178 828 -2160
rect 855 -2178 864 -2160
rect 882 -2178 900 -2151
rect 927 -2178 936 -2151
rect 369 -2214 405 -2205
rect 369 -2232 378 -2214
rect 396 -2232 405 -2214
rect 423 -2232 567 -2205
rect 585 -2223 594 -2205
rect 612 -2223 621 -2205
rect 585 -2232 621 -2223
rect 1395 -2151 1431 -2142
rect 1395 -2169 1404 -2151
rect 1422 -2169 1431 -2151
rect 1449 -2169 1593 -2142
rect 1611 -2160 1620 -2142
rect 1638 -2160 1647 -2142
rect 1611 -2169 1647 -2160
rect 1845 -2097 1890 -2088
rect 1845 -2115 1854 -2097
rect 1881 -2115 1890 -2097
rect 1908 -2115 1926 -2088
rect 1953 -2115 1962 -2088
rect 1044 -2574 1053 -2556
rect 1071 -2574 1080 -2556
rect 1044 -2583 1080 -2574
rect 1098 -2574 1107 -2556
rect 1098 -2583 1125 -2574
rect 1134 -2574 1143 -2556
rect 1161 -2574 1170 -2556
rect 1134 -2583 1170 -2574
rect 1188 -2574 1197 -2556
rect 1188 -2583 1215 -2574
rect 1260 -2574 1269 -2556
rect 1287 -2574 1296 -2556
rect 1260 -2583 1296 -2574
rect 1314 -2574 1323 -2556
rect 1341 -2574 1350 -2556
rect 1314 -2583 1350 -2574
rect 252 -3168 306 -3159
rect 252 -3204 261 -3168
rect 297 -3204 306 -3168
rect 252 -3213 306 -3204
rect 252 -3240 306 -3231
rect 252 -3276 261 -3240
rect 297 -3276 306 -3240
rect 252 -3285 306 -3276
rect 252 -3339 306 -3330
rect 252 -3375 261 -3339
rect 297 -3375 306 -3339
rect 252 -3384 306 -3375
rect 1062 -3168 1116 -3159
rect 1062 -3204 1071 -3168
rect 1107 -3204 1116 -3168
rect 1062 -3213 1116 -3204
rect 252 -3411 306 -3402
rect 252 -3447 261 -3411
rect 297 -3447 306 -3411
rect 252 -3456 306 -3447
rect 252 -3528 306 -3519
rect 252 -3564 261 -3528
rect 297 -3564 306 -3528
rect 252 -3582 306 -3564
rect 252 -3609 306 -3600
rect 252 -3645 261 -3609
rect 297 -3645 306 -3609
rect 252 -3654 306 -3645
rect 252 -3690 306 -3681
rect 252 -3726 261 -3690
rect 297 -3726 306 -3690
rect 252 -3744 306 -3726
rect 252 -3771 306 -3762
rect 252 -3807 261 -3771
rect 297 -3807 306 -3771
rect 252 -3816 306 -3807
rect 1062 -3240 1116 -3231
rect 1062 -3276 1071 -3240
rect 1107 -3276 1116 -3240
rect 1062 -3285 1116 -3276
rect 1062 -3339 1116 -3330
rect 1062 -3375 1071 -3339
rect 1107 -3375 1116 -3339
rect 1062 -3384 1116 -3375
rect 1944 -3168 1998 -3159
rect 1944 -3204 1953 -3168
rect 1989 -3204 1998 -3168
rect 1944 -3213 1998 -3204
rect 1062 -3411 1116 -3402
rect 1062 -3447 1071 -3411
rect 1107 -3447 1116 -3411
rect 1062 -3456 1116 -3447
rect 1062 -3528 1116 -3519
rect 1062 -3564 1071 -3528
rect 1107 -3564 1116 -3528
rect 1062 -3582 1116 -3564
rect 1062 -3609 1116 -3600
rect 1062 -3645 1071 -3609
rect 1107 -3645 1116 -3609
rect 1062 -3654 1116 -3645
rect 1062 -3690 1116 -3681
rect 1062 -3726 1071 -3690
rect 1107 -3726 1116 -3690
rect 1062 -3744 1116 -3726
rect 1062 -3771 1116 -3762
rect 1062 -3807 1071 -3771
rect 1107 -3807 1116 -3771
rect 1062 -3816 1116 -3807
rect 1944 -3240 1998 -3231
rect 1944 -3276 1953 -3240
rect 1989 -3276 1998 -3240
rect 1944 -3285 1998 -3276
rect 1944 -3339 1998 -3330
rect 1944 -3375 1953 -3339
rect 1989 -3375 1998 -3339
rect 1944 -3384 1998 -3375
rect 1944 -3411 1998 -3402
rect 1944 -3447 1953 -3411
rect 1989 -3447 1998 -3411
rect 1944 -3456 1998 -3447
rect 1944 -3528 1998 -3519
rect 1944 -3564 1953 -3528
rect 1989 -3564 1998 -3528
rect 1944 -3582 1998 -3564
rect 1944 -3609 1998 -3600
rect 1944 -3645 1953 -3609
rect 1989 -3645 1998 -3609
rect 1944 -3654 1998 -3645
rect 1944 -3690 1998 -3681
rect 1944 -3726 1953 -3690
rect 1989 -3726 1998 -3690
rect 1944 -3744 1998 -3726
rect 1944 -3771 1998 -3762
rect 1944 -3807 1953 -3771
rect 1989 -3807 1998 -3771
rect 1944 -3816 1998 -3807
rect 819 -4257 864 -4248
rect 819 -4275 828 -4257
rect 855 -4275 864 -4257
rect 882 -4275 900 -4248
rect 927 -4275 936 -4248
rect 369 -4311 405 -4302
rect 369 -4329 378 -4311
rect 396 -4329 405 -4311
rect 423 -4329 567 -4302
rect 585 -4320 594 -4302
rect 612 -4320 621 -4302
rect 585 -4329 621 -4320
rect 1395 -4248 1431 -4239
rect 1395 -4266 1404 -4248
rect 1422 -4266 1431 -4248
rect 1449 -4266 1593 -4239
rect 1611 -4257 1620 -4239
rect 1638 -4257 1647 -4239
rect 1611 -4266 1647 -4257
rect 1845 -4194 1890 -4185
rect 1845 -4212 1854 -4194
rect 1881 -4212 1890 -4194
rect 1908 -4212 1926 -4185
rect 1953 -4212 1962 -4185
rect 1044 -4671 1053 -4653
rect 1071 -4671 1080 -4653
rect 1044 -4680 1080 -4671
rect 1098 -4671 1107 -4653
rect 1098 -4680 1125 -4671
rect 1134 -4671 1143 -4653
rect 1161 -4671 1170 -4653
rect 1134 -4680 1170 -4671
rect 1188 -4671 1197 -4653
rect 1188 -4680 1215 -4671
rect 1260 -4671 1269 -4653
rect 1287 -4671 1296 -4653
rect 1260 -4680 1296 -4671
rect 1314 -4671 1323 -4653
rect 1341 -4671 1350 -4653
rect 1314 -4680 1350 -4671
rect 252 -5283 306 -5274
rect 252 -5319 261 -5283
rect 297 -5319 306 -5283
rect 252 -5328 306 -5319
rect 252 -5355 306 -5346
rect 252 -5391 261 -5355
rect 297 -5391 306 -5355
rect 252 -5400 306 -5391
rect 252 -5454 306 -5445
rect 252 -5490 261 -5454
rect 297 -5490 306 -5454
rect 252 -5499 306 -5490
rect 1062 -5283 1116 -5274
rect 1062 -5319 1071 -5283
rect 1107 -5319 1116 -5283
rect 1062 -5328 1116 -5319
rect 252 -5526 306 -5517
rect 252 -5562 261 -5526
rect 297 -5562 306 -5526
rect 252 -5571 306 -5562
rect 252 -5643 306 -5634
rect 252 -5679 261 -5643
rect 297 -5679 306 -5643
rect 252 -5697 306 -5679
rect 252 -5724 306 -5715
rect 252 -5760 261 -5724
rect 297 -5760 306 -5724
rect 252 -5769 306 -5760
rect 252 -5805 306 -5796
rect 252 -5841 261 -5805
rect 297 -5841 306 -5805
rect 252 -5859 306 -5841
rect 252 -5886 306 -5877
rect 252 -5922 261 -5886
rect 297 -5922 306 -5886
rect 252 -5931 306 -5922
rect 1062 -5355 1116 -5346
rect 1062 -5391 1071 -5355
rect 1107 -5391 1116 -5355
rect 1062 -5400 1116 -5391
rect 1062 -5454 1116 -5445
rect 1062 -5490 1071 -5454
rect 1107 -5490 1116 -5454
rect 1062 -5499 1116 -5490
rect 1944 -5283 1998 -5274
rect 1944 -5319 1953 -5283
rect 1989 -5319 1998 -5283
rect 1944 -5328 1998 -5319
rect 1062 -5526 1116 -5517
rect 1062 -5562 1071 -5526
rect 1107 -5562 1116 -5526
rect 1062 -5571 1116 -5562
rect 1062 -5643 1116 -5634
rect 1062 -5679 1071 -5643
rect 1107 -5679 1116 -5643
rect 1062 -5697 1116 -5679
rect 1062 -5724 1116 -5715
rect 1062 -5760 1071 -5724
rect 1107 -5760 1116 -5724
rect 1062 -5769 1116 -5760
rect 1062 -5805 1116 -5796
rect 1062 -5841 1071 -5805
rect 1107 -5841 1116 -5805
rect 1062 -5859 1116 -5841
rect 1062 -5886 1116 -5877
rect 1062 -5922 1071 -5886
rect 1107 -5922 1116 -5886
rect 1062 -5931 1116 -5922
rect 1944 -5355 1998 -5346
rect 1944 -5391 1953 -5355
rect 1989 -5391 1998 -5355
rect 1944 -5400 1998 -5391
rect 1944 -5454 1998 -5445
rect 1944 -5490 1953 -5454
rect 1989 -5490 1998 -5454
rect 1944 -5499 1998 -5490
rect 1944 -5526 1998 -5517
rect 1944 -5562 1953 -5526
rect 1989 -5562 1998 -5526
rect 1944 -5571 1998 -5562
rect 1944 -5643 1998 -5634
rect 1944 -5679 1953 -5643
rect 1989 -5679 1998 -5643
rect 1944 -5697 1998 -5679
rect 1944 -5724 1998 -5715
rect 1944 -5760 1953 -5724
rect 1989 -5760 1998 -5724
rect 1944 -5769 1998 -5760
rect 1944 -5805 1998 -5796
rect 1944 -5841 1953 -5805
rect 1989 -5841 1998 -5805
rect 1944 -5859 1998 -5841
rect 1944 -5886 1998 -5877
rect 1944 -5922 1953 -5886
rect 1989 -5922 1998 -5886
rect 1944 -5931 1998 -5922
rect 819 -6372 864 -6363
rect 819 -6390 828 -6372
rect 855 -6390 864 -6372
rect 882 -6390 900 -6363
rect 927 -6390 936 -6363
rect 369 -6426 405 -6417
rect 369 -6444 378 -6426
rect 396 -6444 405 -6426
rect 423 -6444 567 -6417
rect 585 -6435 594 -6417
rect 612 -6435 621 -6417
rect 585 -6444 621 -6435
rect 1395 -6363 1431 -6354
rect 1395 -6381 1404 -6363
rect 1422 -6381 1431 -6363
rect 1449 -6381 1593 -6354
rect 1611 -6372 1620 -6354
rect 1638 -6372 1647 -6354
rect 1611 -6381 1647 -6372
rect 1845 -6309 1890 -6300
rect 1845 -6327 1854 -6309
rect 1881 -6327 1890 -6309
rect 1908 -6327 1926 -6300
rect 1953 -6327 1962 -6300
rect 1044 -6786 1053 -6768
rect 1071 -6786 1080 -6768
rect 1044 -6795 1080 -6786
rect 1098 -6786 1107 -6768
rect 1098 -6795 1125 -6786
rect 1134 -6786 1143 -6768
rect 1161 -6786 1170 -6768
rect 1134 -6795 1170 -6786
rect 1188 -6786 1197 -6768
rect 1188 -6795 1215 -6786
rect 1260 -6786 1269 -6768
rect 1287 -6786 1296 -6768
rect 1260 -6795 1296 -6786
rect 1314 -6786 1323 -6768
rect 1341 -6786 1350 -6768
rect 1314 -6795 1350 -6786
rect 252 -7218 306 -7209
rect 252 -7254 261 -7218
rect 297 -7254 306 -7218
rect 252 -7263 306 -7254
rect 252 -7290 306 -7281
rect 252 -7326 261 -7290
rect 297 -7326 306 -7290
rect 252 -7335 306 -7326
rect 252 -7389 306 -7380
rect 252 -7425 261 -7389
rect 297 -7425 306 -7389
rect 252 -7434 306 -7425
rect 1062 -7218 1116 -7209
rect 1062 -7254 1071 -7218
rect 1107 -7254 1116 -7218
rect 1062 -7263 1116 -7254
rect 252 -7461 306 -7452
rect 252 -7497 261 -7461
rect 297 -7497 306 -7461
rect 252 -7506 306 -7497
rect 252 -7578 306 -7569
rect 252 -7614 261 -7578
rect 297 -7614 306 -7578
rect 252 -7632 306 -7614
rect 252 -7659 306 -7650
rect 252 -7695 261 -7659
rect 297 -7695 306 -7659
rect 252 -7704 306 -7695
rect 252 -7740 306 -7731
rect 252 -7776 261 -7740
rect 297 -7776 306 -7740
rect 252 -7794 306 -7776
rect 252 -7821 306 -7812
rect 252 -7857 261 -7821
rect 297 -7857 306 -7821
rect 252 -7866 306 -7857
rect 1062 -7290 1116 -7281
rect 1062 -7326 1071 -7290
rect 1107 -7326 1116 -7290
rect 1062 -7335 1116 -7326
rect 1062 -7389 1116 -7380
rect 1062 -7425 1071 -7389
rect 1107 -7425 1116 -7389
rect 1062 -7434 1116 -7425
rect 1944 -7218 1998 -7209
rect 1944 -7254 1953 -7218
rect 1989 -7254 1998 -7218
rect 1944 -7263 1998 -7254
rect 1062 -7461 1116 -7452
rect 1062 -7497 1071 -7461
rect 1107 -7497 1116 -7461
rect 1062 -7506 1116 -7497
rect 1062 -7578 1116 -7569
rect 1062 -7614 1071 -7578
rect 1107 -7614 1116 -7578
rect 1062 -7632 1116 -7614
rect 1062 -7659 1116 -7650
rect 1062 -7695 1071 -7659
rect 1107 -7695 1116 -7659
rect 1062 -7704 1116 -7695
rect 1062 -7740 1116 -7731
rect 1062 -7776 1071 -7740
rect 1107 -7776 1116 -7740
rect 1062 -7794 1116 -7776
rect 1062 -7821 1116 -7812
rect 1062 -7857 1071 -7821
rect 1107 -7857 1116 -7821
rect 1062 -7866 1116 -7857
rect 1944 -7290 1998 -7281
rect 1944 -7326 1953 -7290
rect 1989 -7326 1998 -7290
rect 1944 -7335 1998 -7326
rect 1944 -7389 1998 -7380
rect 1944 -7425 1953 -7389
rect 1989 -7425 1998 -7389
rect 1944 -7434 1998 -7425
rect 1944 -7461 1998 -7452
rect 1944 -7497 1953 -7461
rect 1989 -7497 1998 -7461
rect 1944 -7506 1998 -7497
rect 1944 -7578 1998 -7569
rect 1944 -7614 1953 -7578
rect 1989 -7614 1998 -7578
rect 1944 -7632 1998 -7614
rect 1944 -7659 1998 -7650
rect 1944 -7695 1953 -7659
rect 1989 -7695 1998 -7659
rect 1944 -7704 1998 -7695
rect 1944 -7740 1998 -7731
rect 1944 -7776 1953 -7740
rect 1989 -7776 1998 -7740
rect 1944 -7794 1998 -7776
rect 1944 -7821 1998 -7812
rect 1944 -7857 1953 -7821
rect 1989 -7857 1998 -7821
rect 1944 -7866 1998 -7857
rect 819 -8307 864 -8298
rect 819 -8325 828 -8307
rect 855 -8325 864 -8307
rect 882 -8325 900 -8298
rect 927 -8325 936 -8298
rect 369 -8361 405 -8352
rect 369 -8379 378 -8361
rect 396 -8379 405 -8361
rect 423 -8379 567 -8352
rect 585 -8370 594 -8352
rect 612 -8370 621 -8352
rect 585 -8379 621 -8370
rect 1395 -8298 1431 -8289
rect 1395 -8316 1404 -8298
rect 1422 -8316 1431 -8298
rect 1449 -8316 1593 -8289
rect 1611 -8307 1620 -8289
rect 1638 -8307 1647 -8289
rect 1611 -8316 1647 -8307
rect 1845 -8244 1890 -8235
rect 1845 -8262 1854 -8244
rect 1881 -8262 1890 -8244
rect 1908 -8262 1926 -8235
rect 1953 -8262 1962 -8235
rect 1044 -8721 1053 -8703
rect 1071 -8721 1080 -8703
rect 1044 -8730 1080 -8721
rect 1098 -8721 1107 -8703
rect 1098 -8730 1125 -8721
rect 1134 -8721 1143 -8703
rect 1161 -8721 1170 -8703
rect 1134 -8730 1170 -8721
rect 1188 -8721 1197 -8703
rect 1188 -8730 1215 -8721
rect 1260 -8721 1269 -8703
rect 1287 -8721 1296 -8703
rect 1260 -8730 1296 -8721
rect 1314 -8721 1323 -8703
rect 1341 -8721 1350 -8703
rect 1314 -8730 1350 -8721
<< pdiffusion >>
rect 504 -1071 567 -1062
rect 504 -1107 513 -1071
rect 549 -1107 567 -1071
rect 504 -1116 567 -1107
rect 504 -1143 567 -1134
rect 504 -1179 513 -1143
rect 549 -1179 567 -1143
rect 504 -1188 567 -1179
rect 504 -1242 567 -1233
rect 504 -1278 513 -1242
rect 549 -1278 567 -1242
rect 504 -1287 567 -1278
rect 1314 -1071 1377 -1062
rect 1314 -1107 1323 -1071
rect 1359 -1107 1377 -1071
rect 1314 -1116 1377 -1107
rect 504 -1314 567 -1305
rect 504 -1350 513 -1314
rect 549 -1350 567 -1314
rect 504 -1359 567 -1350
rect 504 -1431 567 -1422
rect 504 -1467 513 -1431
rect 549 -1467 567 -1431
rect 504 -1485 567 -1467
rect 504 -1512 567 -1503
rect 504 -1548 513 -1512
rect 549 -1548 567 -1512
rect 504 -1557 567 -1548
rect 504 -1593 567 -1584
rect 504 -1629 513 -1593
rect 549 -1629 567 -1593
rect 504 -1647 567 -1629
rect 504 -1674 567 -1665
rect 504 -1710 513 -1674
rect 549 -1710 567 -1674
rect 504 -1719 567 -1710
rect 1314 -1143 1377 -1134
rect 1314 -1179 1323 -1143
rect 1359 -1179 1377 -1143
rect 1314 -1188 1377 -1179
rect 1314 -1242 1377 -1233
rect 1314 -1278 1323 -1242
rect 1359 -1278 1377 -1242
rect 1314 -1287 1377 -1278
rect 2196 -1071 2259 -1062
rect 2196 -1107 2205 -1071
rect 2241 -1107 2259 -1071
rect 2196 -1116 2259 -1107
rect 1314 -1314 1377 -1305
rect 1314 -1350 1323 -1314
rect 1359 -1350 1377 -1314
rect 1314 -1359 1377 -1350
rect 1314 -1431 1377 -1422
rect 1314 -1467 1323 -1431
rect 1359 -1467 1377 -1431
rect 1314 -1485 1377 -1467
rect 1314 -1512 1377 -1503
rect 1314 -1548 1323 -1512
rect 1359 -1548 1377 -1512
rect 1314 -1557 1377 -1548
rect 1314 -1593 1377 -1584
rect 1314 -1629 1323 -1593
rect 1359 -1629 1377 -1593
rect 1314 -1647 1377 -1629
rect 1314 -1674 1377 -1665
rect 1314 -1710 1323 -1674
rect 1359 -1710 1377 -1674
rect 1314 -1719 1377 -1710
rect 2196 -1143 2259 -1134
rect 2196 -1179 2205 -1143
rect 2241 -1179 2259 -1143
rect 2196 -1188 2259 -1179
rect 2196 -1242 2259 -1233
rect 2196 -1278 2205 -1242
rect 2241 -1278 2259 -1242
rect 2196 -1287 2259 -1278
rect 2196 -1314 2259 -1305
rect 2196 -1350 2205 -1314
rect 2241 -1350 2259 -1314
rect 2196 -1359 2259 -1350
rect 2196 -1431 2259 -1422
rect 2196 -1467 2205 -1431
rect 2241 -1467 2259 -1431
rect 2196 -1485 2259 -1467
rect 2196 -1512 2259 -1503
rect 2196 -1548 2205 -1512
rect 2241 -1548 2259 -1512
rect 2196 -1557 2259 -1548
rect 2196 -1593 2259 -1584
rect 2196 -1629 2205 -1593
rect 2241 -1629 2259 -1593
rect 2196 -1647 2259 -1629
rect 2196 -1674 2259 -1665
rect 2196 -1710 2205 -1674
rect 2241 -1710 2259 -1674
rect 2196 -1719 2259 -1710
rect 369 -2070 405 -2061
rect 369 -2088 378 -2070
rect 396 -2088 405 -2070
rect 369 -2106 405 -2088
rect 423 -2079 486 -2061
rect 423 -2097 432 -2079
rect 450 -2097 486 -2079
rect 423 -2106 486 -2097
rect 522 -2070 567 -2061
rect 522 -2088 531 -2070
rect 549 -2088 567 -2070
rect 522 -2106 567 -2088
rect 585 -2070 621 -2061
rect 585 -2088 594 -2070
rect 612 -2088 621 -2070
rect 585 -2106 621 -2088
rect 819 -2052 828 -2025
rect 855 -2052 864 -2025
rect 819 -2079 864 -2052
rect 882 -2034 936 -2025
rect 882 -2061 900 -2034
rect 927 -2061 936 -2034
rect 882 -2079 936 -2061
rect 1395 -2007 1431 -1998
rect 1395 -2025 1404 -2007
rect 1422 -2025 1431 -2007
rect 1395 -2043 1431 -2025
rect 1449 -2016 1512 -1998
rect 1449 -2034 1458 -2016
rect 1476 -2034 1512 -2016
rect 1449 -2043 1512 -2034
rect 1548 -2007 1593 -1998
rect 1548 -2025 1557 -2007
rect 1575 -2025 1593 -2007
rect 1548 -2043 1593 -2025
rect 1611 -2007 1647 -1998
rect 1611 -2025 1620 -2007
rect 1638 -2025 1647 -2007
rect 1611 -2043 1647 -2025
rect 1845 -1989 1854 -1962
rect 1881 -1989 1890 -1962
rect 1845 -2016 1890 -1989
rect 1908 -1971 1962 -1962
rect 1908 -1998 1926 -1971
rect 1953 -1998 1962 -1971
rect 1908 -2016 1962 -1998
rect 1035 -2430 1080 -2421
rect 1035 -2448 1044 -2430
rect 1062 -2448 1080 -2430
rect 1035 -2466 1080 -2448
rect 1098 -2466 1170 -2421
rect 1188 -2439 1215 -2421
rect 1188 -2457 1197 -2439
rect 1188 -2466 1215 -2457
rect 1260 -2430 1296 -2421
rect 1260 -2448 1269 -2430
rect 1287 -2448 1296 -2430
rect 1260 -2466 1296 -2448
rect 1314 -2439 1350 -2421
rect 1314 -2457 1323 -2439
rect 1341 -2457 1350 -2439
rect 1314 -2466 1350 -2457
rect 504 -3168 567 -3159
rect 504 -3204 513 -3168
rect 549 -3204 567 -3168
rect 504 -3213 567 -3204
rect 504 -3240 567 -3231
rect 504 -3276 513 -3240
rect 549 -3276 567 -3240
rect 504 -3285 567 -3276
rect 504 -3339 567 -3330
rect 504 -3375 513 -3339
rect 549 -3375 567 -3339
rect 504 -3384 567 -3375
rect 1314 -3168 1377 -3159
rect 1314 -3204 1323 -3168
rect 1359 -3204 1377 -3168
rect 1314 -3213 1377 -3204
rect 504 -3411 567 -3402
rect 504 -3447 513 -3411
rect 549 -3447 567 -3411
rect 504 -3456 567 -3447
rect 504 -3528 567 -3519
rect 504 -3564 513 -3528
rect 549 -3564 567 -3528
rect 504 -3582 567 -3564
rect 504 -3609 567 -3600
rect 504 -3645 513 -3609
rect 549 -3645 567 -3609
rect 504 -3654 567 -3645
rect 504 -3690 567 -3681
rect 504 -3726 513 -3690
rect 549 -3726 567 -3690
rect 504 -3744 567 -3726
rect 504 -3771 567 -3762
rect 504 -3807 513 -3771
rect 549 -3807 567 -3771
rect 504 -3816 567 -3807
rect 1314 -3240 1377 -3231
rect 1314 -3276 1323 -3240
rect 1359 -3276 1377 -3240
rect 1314 -3285 1377 -3276
rect 1314 -3339 1377 -3330
rect 1314 -3375 1323 -3339
rect 1359 -3375 1377 -3339
rect 1314 -3384 1377 -3375
rect 2196 -3168 2259 -3159
rect 2196 -3204 2205 -3168
rect 2241 -3204 2259 -3168
rect 2196 -3213 2259 -3204
rect 1314 -3411 1377 -3402
rect 1314 -3447 1323 -3411
rect 1359 -3447 1377 -3411
rect 1314 -3456 1377 -3447
rect 1314 -3528 1377 -3519
rect 1314 -3564 1323 -3528
rect 1359 -3564 1377 -3528
rect 1314 -3582 1377 -3564
rect 1314 -3609 1377 -3600
rect 1314 -3645 1323 -3609
rect 1359 -3645 1377 -3609
rect 1314 -3654 1377 -3645
rect 1314 -3690 1377 -3681
rect 1314 -3726 1323 -3690
rect 1359 -3726 1377 -3690
rect 1314 -3744 1377 -3726
rect 1314 -3771 1377 -3762
rect 1314 -3807 1323 -3771
rect 1359 -3807 1377 -3771
rect 1314 -3816 1377 -3807
rect 2196 -3240 2259 -3231
rect 2196 -3276 2205 -3240
rect 2241 -3276 2259 -3240
rect 2196 -3285 2259 -3276
rect 2196 -3339 2259 -3330
rect 2196 -3375 2205 -3339
rect 2241 -3375 2259 -3339
rect 2196 -3384 2259 -3375
rect 2196 -3411 2259 -3402
rect 2196 -3447 2205 -3411
rect 2241 -3447 2259 -3411
rect 2196 -3456 2259 -3447
rect 2196 -3528 2259 -3519
rect 2196 -3564 2205 -3528
rect 2241 -3564 2259 -3528
rect 2196 -3582 2259 -3564
rect 2196 -3609 2259 -3600
rect 2196 -3645 2205 -3609
rect 2241 -3645 2259 -3609
rect 2196 -3654 2259 -3645
rect 2196 -3690 2259 -3681
rect 2196 -3726 2205 -3690
rect 2241 -3726 2259 -3690
rect 2196 -3744 2259 -3726
rect 2196 -3771 2259 -3762
rect 2196 -3807 2205 -3771
rect 2241 -3807 2259 -3771
rect 2196 -3816 2259 -3807
rect 369 -4167 405 -4158
rect 369 -4185 378 -4167
rect 396 -4185 405 -4167
rect 369 -4203 405 -4185
rect 423 -4176 486 -4158
rect 423 -4194 432 -4176
rect 450 -4194 486 -4176
rect 423 -4203 486 -4194
rect 522 -4167 567 -4158
rect 522 -4185 531 -4167
rect 549 -4185 567 -4167
rect 522 -4203 567 -4185
rect 585 -4167 621 -4158
rect 585 -4185 594 -4167
rect 612 -4185 621 -4167
rect 585 -4203 621 -4185
rect 819 -4149 828 -4122
rect 855 -4149 864 -4122
rect 819 -4176 864 -4149
rect 882 -4131 936 -4122
rect 882 -4158 900 -4131
rect 927 -4158 936 -4131
rect 882 -4176 936 -4158
rect 1395 -4104 1431 -4095
rect 1395 -4122 1404 -4104
rect 1422 -4122 1431 -4104
rect 1395 -4140 1431 -4122
rect 1449 -4113 1512 -4095
rect 1449 -4131 1458 -4113
rect 1476 -4131 1512 -4113
rect 1449 -4140 1512 -4131
rect 1548 -4104 1593 -4095
rect 1548 -4122 1557 -4104
rect 1575 -4122 1593 -4104
rect 1548 -4140 1593 -4122
rect 1611 -4104 1647 -4095
rect 1611 -4122 1620 -4104
rect 1638 -4122 1647 -4104
rect 1611 -4140 1647 -4122
rect 1845 -4086 1854 -4059
rect 1881 -4086 1890 -4059
rect 1845 -4113 1890 -4086
rect 1908 -4068 1962 -4059
rect 1908 -4095 1926 -4068
rect 1953 -4095 1962 -4068
rect 1908 -4113 1962 -4095
rect 1035 -4527 1080 -4518
rect 1035 -4545 1044 -4527
rect 1062 -4545 1080 -4527
rect 1035 -4563 1080 -4545
rect 1098 -4563 1170 -4518
rect 1188 -4536 1215 -4518
rect 1188 -4554 1197 -4536
rect 1188 -4563 1215 -4554
rect 1260 -4527 1296 -4518
rect 1260 -4545 1269 -4527
rect 1287 -4545 1296 -4527
rect 1260 -4563 1296 -4545
rect 1314 -4536 1350 -4518
rect 1314 -4554 1323 -4536
rect 1341 -4554 1350 -4536
rect 1314 -4563 1350 -4554
rect 504 -5283 567 -5274
rect 504 -5319 513 -5283
rect 549 -5319 567 -5283
rect 504 -5328 567 -5319
rect 504 -5355 567 -5346
rect 504 -5391 513 -5355
rect 549 -5391 567 -5355
rect 504 -5400 567 -5391
rect 504 -5454 567 -5445
rect 504 -5490 513 -5454
rect 549 -5490 567 -5454
rect 504 -5499 567 -5490
rect 1314 -5283 1377 -5274
rect 1314 -5319 1323 -5283
rect 1359 -5319 1377 -5283
rect 1314 -5328 1377 -5319
rect 504 -5526 567 -5517
rect 504 -5562 513 -5526
rect 549 -5562 567 -5526
rect 504 -5571 567 -5562
rect 504 -5643 567 -5634
rect 504 -5679 513 -5643
rect 549 -5679 567 -5643
rect 504 -5697 567 -5679
rect 504 -5724 567 -5715
rect 504 -5760 513 -5724
rect 549 -5760 567 -5724
rect 504 -5769 567 -5760
rect 504 -5805 567 -5796
rect 504 -5841 513 -5805
rect 549 -5841 567 -5805
rect 504 -5859 567 -5841
rect 504 -5886 567 -5877
rect 504 -5922 513 -5886
rect 549 -5922 567 -5886
rect 504 -5931 567 -5922
rect 1314 -5355 1377 -5346
rect 1314 -5391 1323 -5355
rect 1359 -5391 1377 -5355
rect 1314 -5400 1377 -5391
rect 1314 -5454 1377 -5445
rect 1314 -5490 1323 -5454
rect 1359 -5490 1377 -5454
rect 1314 -5499 1377 -5490
rect 2196 -5283 2259 -5274
rect 2196 -5319 2205 -5283
rect 2241 -5319 2259 -5283
rect 2196 -5328 2259 -5319
rect 1314 -5526 1377 -5517
rect 1314 -5562 1323 -5526
rect 1359 -5562 1377 -5526
rect 1314 -5571 1377 -5562
rect 1314 -5643 1377 -5634
rect 1314 -5679 1323 -5643
rect 1359 -5679 1377 -5643
rect 1314 -5697 1377 -5679
rect 1314 -5724 1377 -5715
rect 1314 -5760 1323 -5724
rect 1359 -5760 1377 -5724
rect 1314 -5769 1377 -5760
rect 1314 -5805 1377 -5796
rect 1314 -5841 1323 -5805
rect 1359 -5841 1377 -5805
rect 1314 -5859 1377 -5841
rect 1314 -5886 1377 -5877
rect 1314 -5922 1323 -5886
rect 1359 -5922 1377 -5886
rect 1314 -5931 1377 -5922
rect 2196 -5355 2259 -5346
rect 2196 -5391 2205 -5355
rect 2241 -5391 2259 -5355
rect 2196 -5400 2259 -5391
rect 2196 -5454 2259 -5445
rect 2196 -5490 2205 -5454
rect 2241 -5490 2259 -5454
rect 2196 -5499 2259 -5490
rect 2196 -5526 2259 -5517
rect 2196 -5562 2205 -5526
rect 2241 -5562 2259 -5526
rect 2196 -5571 2259 -5562
rect 2196 -5643 2259 -5634
rect 2196 -5679 2205 -5643
rect 2241 -5679 2259 -5643
rect 2196 -5697 2259 -5679
rect 2196 -5724 2259 -5715
rect 2196 -5760 2205 -5724
rect 2241 -5760 2259 -5724
rect 2196 -5769 2259 -5760
rect 2196 -5805 2259 -5796
rect 2196 -5841 2205 -5805
rect 2241 -5841 2259 -5805
rect 2196 -5859 2259 -5841
rect 2196 -5886 2259 -5877
rect 2196 -5922 2205 -5886
rect 2241 -5922 2259 -5886
rect 2196 -5931 2259 -5922
rect 369 -6282 405 -6273
rect 369 -6300 378 -6282
rect 396 -6300 405 -6282
rect 369 -6318 405 -6300
rect 423 -6291 486 -6273
rect 423 -6309 432 -6291
rect 450 -6309 486 -6291
rect 423 -6318 486 -6309
rect 522 -6282 567 -6273
rect 522 -6300 531 -6282
rect 549 -6300 567 -6282
rect 522 -6318 567 -6300
rect 585 -6282 621 -6273
rect 585 -6300 594 -6282
rect 612 -6300 621 -6282
rect 585 -6318 621 -6300
rect 819 -6264 828 -6237
rect 855 -6264 864 -6237
rect 819 -6291 864 -6264
rect 882 -6246 936 -6237
rect 882 -6273 900 -6246
rect 927 -6273 936 -6246
rect 882 -6291 936 -6273
rect 1395 -6219 1431 -6210
rect 1395 -6237 1404 -6219
rect 1422 -6237 1431 -6219
rect 1395 -6255 1431 -6237
rect 1449 -6228 1512 -6210
rect 1449 -6246 1458 -6228
rect 1476 -6246 1512 -6228
rect 1449 -6255 1512 -6246
rect 1548 -6219 1593 -6210
rect 1548 -6237 1557 -6219
rect 1575 -6237 1593 -6219
rect 1548 -6255 1593 -6237
rect 1611 -6219 1647 -6210
rect 1611 -6237 1620 -6219
rect 1638 -6237 1647 -6219
rect 1611 -6255 1647 -6237
rect 1845 -6201 1854 -6174
rect 1881 -6201 1890 -6174
rect 1845 -6228 1890 -6201
rect 1908 -6183 1962 -6174
rect 1908 -6210 1926 -6183
rect 1953 -6210 1962 -6183
rect 1908 -6228 1962 -6210
rect 1035 -6642 1080 -6633
rect 1035 -6660 1044 -6642
rect 1062 -6660 1080 -6642
rect 1035 -6678 1080 -6660
rect 1098 -6678 1170 -6633
rect 1188 -6651 1215 -6633
rect 1188 -6669 1197 -6651
rect 1188 -6678 1215 -6669
rect 1260 -6642 1296 -6633
rect 1260 -6660 1269 -6642
rect 1287 -6660 1296 -6642
rect 1260 -6678 1296 -6660
rect 1314 -6651 1350 -6633
rect 1314 -6669 1323 -6651
rect 1341 -6669 1350 -6651
rect 1314 -6678 1350 -6669
rect 504 -7218 567 -7209
rect 504 -7254 513 -7218
rect 549 -7254 567 -7218
rect 504 -7263 567 -7254
rect 504 -7290 567 -7281
rect 504 -7326 513 -7290
rect 549 -7326 567 -7290
rect 504 -7335 567 -7326
rect 504 -7389 567 -7380
rect 504 -7425 513 -7389
rect 549 -7425 567 -7389
rect 504 -7434 567 -7425
rect 1314 -7218 1377 -7209
rect 1314 -7254 1323 -7218
rect 1359 -7254 1377 -7218
rect 1314 -7263 1377 -7254
rect 504 -7461 567 -7452
rect 504 -7497 513 -7461
rect 549 -7497 567 -7461
rect 504 -7506 567 -7497
rect 504 -7578 567 -7569
rect 504 -7614 513 -7578
rect 549 -7614 567 -7578
rect 504 -7632 567 -7614
rect 504 -7659 567 -7650
rect 504 -7695 513 -7659
rect 549 -7695 567 -7659
rect 504 -7704 567 -7695
rect 504 -7740 567 -7731
rect 504 -7776 513 -7740
rect 549 -7776 567 -7740
rect 504 -7794 567 -7776
rect 504 -7821 567 -7812
rect 504 -7857 513 -7821
rect 549 -7857 567 -7821
rect 504 -7866 567 -7857
rect 1314 -7290 1377 -7281
rect 1314 -7326 1323 -7290
rect 1359 -7326 1377 -7290
rect 1314 -7335 1377 -7326
rect 1314 -7389 1377 -7380
rect 1314 -7425 1323 -7389
rect 1359 -7425 1377 -7389
rect 1314 -7434 1377 -7425
rect 2196 -7218 2259 -7209
rect 2196 -7254 2205 -7218
rect 2241 -7254 2259 -7218
rect 2196 -7263 2259 -7254
rect 1314 -7461 1377 -7452
rect 1314 -7497 1323 -7461
rect 1359 -7497 1377 -7461
rect 1314 -7506 1377 -7497
rect 1314 -7578 1377 -7569
rect 1314 -7614 1323 -7578
rect 1359 -7614 1377 -7578
rect 1314 -7632 1377 -7614
rect 1314 -7659 1377 -7650
rect 1314 -7695 1323 -7659
rect 1359 -7695 1377 -7659
rect 1314 -7704 1377 -7695
rect 1314 -7740 1377 -7731
rect 1314 -7776 1323 -7740
rect 1359 -7776 1377 -7740
rect 1314 -7794 1377 -7776
rect 1314 -7821 1377 -7812
rect 1314 -7857 1323 -7821
rect 1359 -7857 1377 -7821
rect 1314 -7866 1377 -7857
rect 2196 -7290 2259 -7281
rect 2196 -7326 2205 -7290
rect 2241 -7326 2259 -7290
rect 2196 -7335 2259 -7326
rect 2196 -7389 2259 -7380
rect 2196 -7425 2205 -7389
rect 2241 -7425 2259 -7389
rect 2196 -7434 2259 -7425
rect 2196 -7461 2259 -7452
rect 2196 -7497 2205 -7461
rect 2241 -7497 2259 -7461
rect 2196 -7506 2259 -7497
rect 2196 -7578 2259 -7569
rect 2196 -7614 2205 -7578
rect 2241 -7614 2259 -7578
rect 2196 -7632 2259 -7614
rect 2196 -7659 2259 -7650
rect 2196 -7695 2205 -7659
rect 2241 -7695 2259 -7659
rect 2196 -7704 2259 -7695
rect 2196 -7740 2259 -7731
rect 2196 -7776 2205 -7740
rect 2241 -7776 2259 -7740
rect 2196 -7794 2259 -7776
rect 2196 -7821 2259 -7812
rect 2196 -7857 2205 -7821
rect 2241 -7857 2259 -7821
rect 2196 -7866 2259 -7857
rect 369 -8217 405 -8208
rect 369 -8235 378 -8217
rect 396 -8235 405 -8217
rect 369 -8253 405 -8235
rect 423 -8226 486 -8208
rect 423 -8244 432 -8226
rect 450 -8244 486 -8226
rect 423 -8253 486 -8244
rect 522 -8217 567 -8208
rect 522 -8235 531 -8217
rect 549 -8235 567 -8217
rect 522 -8253 567 -8235
rect 585 -8217 621 -8208
rect 585 -8235 594 -8217
rect 612 -8235 621 -8217
rect 585 -8253 621 -8235
rect 819 -8199 828 -8172
rect 855 -8199 864 -8172
rect 819 -8226 864 -8199
rect 882 -8181 936 -8172
rect 882 -8208 900 -8181
rect 927 -8208 936 -8181
rect 882 -8226 936 -8208
rect 1395 -8154 1431 -8145
rect 1395 -8172 1404 -8154
rect 1422 -8172 1431 -8154
rect 1395 -8190 1431 -8172
rect 1449 -8163 1512 -8145
rect 1449 -8181 1458 -8163
rect 1476 -8181 1512 -8163
rect 1449 -8190 1512 -8181
rect 1548 -8154 1593 -8145
rect 1548 -8172 1557 -8154
rect 1575 -8172 1593 -8154
rect 1548 -8190 1593 -8172
rect 1611 -8154 1647 -8145
rect 1611 -8172 1620 -8154
rect 1638 -8172 1647 -8154
rect 1611 -8190 1647 -8172
rect 1845 -8136 1854 -8109
rect 1881 -8136 1890 -8109
rect 1845 -8163 1890 -8136
rect 1908 -8118 1962 -8109
rect 1908 -8145 1926 -8118
rect 1953 -8145 1962 -8118
rect 1908 -8163 1962 -8145
rect 1035 -8577 1080 -8568
rect 1035 -8595 1044 -8577
rect 1062 -8595 1080 -8577
rect 1035 -8613 1080 -8595
rect 1098 -8613 1170 -8568
rect 1188 -8586 1215 -8568
rect 1188 -8604 1197 -8586
rect 1188 -8613 1215 -8604
rect 1260 -8577 1296 -8568
rect 1260 -8595 1269 -8577
rect 1287 -8595 1296 -8577
rect 1260 -8613 1296 -8595
rect 1314 -8586 1350 -8568
rect 1314 -8604 1323 -8586
rect 1341 -8604 1350 -8586
rect 1314 -8613 1350 -8604
<< ndcontact >>
rect 261 -1107 297 -1071
rect 261 -1179 297 -1143
rect 261 -1278 297 -1242
rect 1071 -1107 1107 -1071
rect 261 -1350 297 -1314
rect 261 -1467 297 -1431
rect 261 -1548 297 -1512
rect 261 -1629 297 -1593
rect 261 -1710 297 -1674
rect 1071 -1179 1107 -1143
rect 1071 -1278 1107 -1242
rect 1953 -1107 1989 -1071
rect 1071 -1350 1107 -1314
rect 1071 -1467 1107 -1431
rect 1071 -1548 1107 -1512
rect 1071 -1629 1107 -1593
rect 1071 -1710 1107 -1674
rect 1953 -1179 1989 -1143
rect 1953 -1278 1989 -1242
rect 1953 -1350 1989 -1314
rect 1953 -1467 1989 -1431
rect 1953 -1548 1989 -1512
rect 1953 -1629 1989 -1593
rect 1953 -1710 1989 -1674
rect 828 -2187 855 -2160
rect 900 -2178 927 -2151
rect 378 -2232 396 -2214
rect 594 -2223 612 -2205
rect 1404 -2169 1422 -2151
rect 1620 -2160 1638 -2142
rect 1854 -2124 1881 -2097
rect 1926 -2115 1953 -2088
rect 1053 -2574 1071 -2556
rect 1107 -2574 1125 -2556
rect 1143 -2574 1161 -2556
rect 1197 -2574 1215 -2556
rect 1269 -2574 1287 -2556
rect 1323 -2574 1341 -2556
rect 261 -3204 297 -3168
rect 261 -3276 297 -3240
rect 261 -3375 297 -3339
rect 1071 -3204 1107 -3168
rect 261 -3447 297 -3411
rect 261 -3564 297 -3528
rect 261 -3645 297 -3609
rect 261 -3726 297 -3690
rect 261 -3807 297 -3771
rect 1071 -3276 1107 -3240
rect 1071 -3375 1107 -3339
rect 1953 -3204 1989 -3168
rect 1071 -3447 1107 -3411
rect 1071 -3564 1107 -3528
rect 1071 -3645 1107 -3609
rect 1071 -3726 1107 -3690
rect 1071 -3807 1107 -3771
rect 1953 -3276 1989 -3240
rect 1953 -3375 1989 -3339
rect 1953 -3447 1989 -3411
rect 1953 -3564 1989 -3528
rect 1953 -3645 1989 -3609
rect 1953 -3726 1989 -3690
rect 1953 -3807 1989 -3771
rect 828 -4284 855 -4257
rect 900 -4275 927 -4248
rect 378 -4329 396 -4311
rect 594 -4320 612 -4302
rect 1404 -4266 1422 -4248
rect 1620 -4257 1638 -4239
rect 1854 -4221 1881 -4194
rect 1926 -4212 1953 -4185
rect 1053 -4671 1071 -4653
rect 1107 -4671 1125 -4653
rect 1143 -4671 1161 -4653
rect 1197 -4671 1215 -4653
rect 1269 -4671 1287 -4653
rect 1323 -4671 1341 -4653
rect 261 -5319 297 -5283
rect 261 -5391 297 -5355
rect 261 -5490 297 -5454
rect 1071 -5319 1107 -5283
rect 261 -5562 297 -5526
rect 261 -5679 297 -5643
rect 261 -5760 297 -5724
rect 261 -5841 297 -5805
rect 261 -5922 297 -5886
rect 1071 -5391 1107 -5355
rect 1071 -5490 1107 -5454
rect 1953 -5319 1989 -5283
rect 1071 -5562 1107 -5526
rect 1071 -5679 1107 -5643
rect 1071 -5760 1107 -5724
rect 1071 -5841 1107 -5805
rect 1071 -5922 1107 -5886
rect 1953 -5391 1989 -5355
rect 1953 -5490 1989 -5454
rect 1953 -5562 1989 -5526
rect 1953 -5679 1989 -5643
rect 1953 -5760 1989 -5724
rect 1953 -5841 1989 -5805
rect 1953 -5922 1989 -5886
rect 828 -6399 855 -6372
rect 900 -6390 927 -6363
rect 378 -6444 396 -6426
rect 594 -6435 612 -6417
rect 1404 -6381 1422 -6363
rect 1620 -6372 1638 -6354
rect 1854 -6336 1881 -6309
rect 1926 -6327 1953 -6300
rect 1053 -6786 1071 -6768
rect 1107 -6786 1125 -6768
rect 1143 -6786 1161 -6768
rect 1197 -6786 1215 -6768
rect 1269 -6786 1287 -6768
rect 1323 -6786 1341 -6768
rect 261 -7254 297 -7218
rect 261 -7326 297 -7290
rect 261 -7425 297 -7389
rect 1071 -7254 1107 -7218
rect 261 -7497 297 -7461
rect 261 -7614 297 -7578
rect 261 -7695 297 -7659
rect 261 -7776 297 -7740
rect 261 -7857 297 -7821
rect 1071 -7326 1107 -7290
rect 1071 -7425 1107 -7389
rect 1953 -7254 1989 -7218
rect 1071 -7497 1107 -7461
rect 1071 -7614 1107 -7578
rect 1071 -7695 1107 -7659
rect 1071 -7776 1107 -7740
rect 1071 -7857 1107 -7821
rect 1953 -7326 1989 -7290
rect 1953 -7425 1989 -7389
rect 1953 -7497 1989 -7461
rect 1953 -7614 1989 -7578
rect 1953 -7695 1989 -7659
rect 1953 -7776 1989 -7740
rect 1953 -7857 1989 -7821
rect 828 -8334 855 -8307
rect 900 -8325 927 -8298
rect 378 -8379 396 -8361
rect 594 -8370 612 -8352
rect 1404 -8316 1422 -8298
rect 1620 -8307 1638 -8289
rect 1854 -8271 1881 -8244
rect 1926 -8262 1953 -8235
rect 1053 -8721 1071 -8703
rect 1107 -8721 1125 -8703
rect 1143 -8721 1161 -8703
rect 1197 -8721 1215 -8703
rect 1269 -8721 1287 -8703
rect 1323 -8721 1341 -8703
<< pdcontact >>
rect 513 -1107 549 -1071
rect 513 -1179 549 -1143
rect 513 -1278 549 -1242
rect 1323 -1107 1359 -1071
rect 513 -1350 549 -1314
rect 513 -1467 549 -1431
rect 513 -1548 549 -1512
rect 513 -1629 549 -1593
rect 513 -1710 549 -1674
rect 1323 -1179 1359 -1143
rect 1323 -1278 1359 -1242
rect 2205 -1107 2241 -1071
rect 1323 -1350 1359 -1314
rect 1323 -1467 1359 -1431
rect 1323 -1548 1359 -1512
rect 1323 -1629 1359 -1593
rect 1323 -1710 1359 -1674
rect 2205 -1179 2241 -1143
rect 2205 -1278 2241 -1242
rect 2205 -1350 2241 -1314
rect 2205 -1467 2241 -1431
rect 2205 -1548 2241 -1512
rect 2205 -1629 2241 -1593
rect 2205 -1710 2241 -1674
rect 378 -2088 396 -2070
rect 432 -2097 450 -2079
rect 531 -2088 549 -2070
rect 594 -2088 612 -2070
rect 828 -2052 855 -2025
rect 900 -2061 927 -2034
rect 1404 -2025 1422 -2007
rect 1458 -2034 1476 -2016
rect 1557 -2025 1575 -2007
rect 1620 -2025 1638 -2007
rect 1854 -1989 1881 -1962
rect 1926 -1998 1953 -1971
rect 1044 -2448 1062 -2430
rect 1197 -2457 1215 -2439
rect 1269 -2448 1287 -2430
rect 1323 -2457 1341 -2439
rect 513 -3204 549 -3168
rect 513 -3276 549 -3240
rect 513 -3375 549 -3339
rect 1323 -3204 1359 -3168
rect 513 -3447 549 -3411
rect 513 -3564 549 -3528
rect 513 -3645 549 -3609
rect 513 -3726 549 -3690
rect 513 -3807 549 -3771
rect 1323 -3276 1359 -3240
rect 1323 -3375 1359 -3339
rect 2205 -3204 2241 -3168
rect 1323 -3447 1359 -3411
rect 1323 -3564 1359 -3528
rect 1323 -3645 1359 -3609
rect 1323 -3726 1359 -3690
rect 1323 -3807 1359 -3771
rect 2205 -3276 2241 -3240
rect 2205 -3375 2241 -3339
rect 2205 -3447 2241 -3411
rect 2205 -3564 2241 -3528
rect 2205 -3645 2241 -3609
rect 2205 -3726 2241 -3690
rect 2205 -3807 2241 -3771
rect 378 -4185 396 -4167
rect 432 -4194 450 -4176
rect 531 -4185 549 -4167
rect 594 -4185 612 -4167
rect 828 -4149 855 -4122
rect 900 -4158 927 -4131
rect 1404 -4122 1422 -4104
rect 1458 -4131 1476 -4113
rect 1557 -4122 1575 -4104
rect 1620 -4122 1638 -4104
rect 1854 -4086 1881 -4059
rect 1926 -4095 1953 -4068
rect 1044 -4545 1062 -4527
rect 1197 -4554 1215 -4536
rect 1269 -4545 1287 -4527
rect 1323 -4554 1341 -4536
rect 513 -5319 549 -5283
rect 513 -5391 549 -5355
rect 513 -5490 549 -5454
rect 1323 -5319 1359 -5283
rect 513 -5562 549 -5526
rect 513 -5679 549 -5643
rect 513 -5760 549 -5724
rect 513 -5841 549 -5805
rect 513 -5922 549 -5886
rect 1323 -5391 1359 -5355
rect 1323 -5490 1359 -5454
rect 2205 -5319 2241 -5283
rect 1323 -5562 1359 -5526
rect 1323 -5679 1359 -5643
rect 1323 -5760 1359 -5724
rect 1323 -5841 1359 -5805
rect 1323 -5922 1359 -5886
rect 2205 -5391 2241 -5355
rect 2205 -5490 2241 -5454
rect 2205 -5562 2241 -5526
rect 2205 -5679 2241 -5643
rect 2205 -5760 2241 -5724
rect 2205 -5841 2241 -5805
rect 2205 -5922 2241 -5886
rect 378 -6300 396 -6282
rect 432 -6309 450 -6291
rect 531 -6300 549 -6282
rect 594 -6300 612 -6282
rect 828 -6264 855 -6237
rect 900 -6273 927 -6246
rect 1404 -6237 1422 -6219
rect 1458 -6246 1476 -6228
rect 1557 -6237 1575 -6219
rect 1620 -6237 1638 -6219
rect 1854 -6201 1881 -6174
rect 1926 -6210 1953 -6183
rect 1044 -6660 1062 -6642
rect 1197 -6669 1215 -6651
rect 1269 -6660 1287 -6642
rect 1323 -6669 1341 -6651
rect 513 -7254 549 -7218
rect 513 -7326 549 -7290
rect 513 -7425 549 -7389
rect 1323 -7254 1359 -7218
rect 513 -7497 549 -7461
rect 513 -7614 549 -7578
rect 513 -7695 549 -7659
rect 513 -7776 549 -7740
rect 513 -7857 549 -7821
rect 1323 -7326 1359 -7290
rect 1323 -7425 1359 -7389
rect 2205 -7254 2241 -7218
rect 1323 -7497 1359 -7461
rect 1323 -7614 1359 -7578
rect 1323 -7695 1359 -7659
rect 1323 -7776 1359 -7740
rect 1323 -7857 1359 -7821
rect 2205 -7326 2241 -7290
rect 2205 -7425 2241 -7389
rect 2205 -7497 2241 -7461
rect 2205 -7614 2241 -7578
rect 2205 -7695 2241 -7659
rect 2205 -7776 2241 -7740
rect 2205 -7857 2241 -7821
rect 378 -8235 396 -8217
rect 432 -8244 450 -8226
rect 531 -8235 549 -8217
rect 594 -8235 612 -8217
rect 828 -8199 855 -8172
rect 900 -8208 927 -8181
rect 1404 -8172 1422 -8154
rect 1458 -8181 1476 -8163
rect 1557 -8172 1575 -8154
rect 1620 -8172 1638 -8154
rect 1854 -8136 1881 -8109
rect 1926 -8145 1953 -8118
rect 1044 -8595 1062 -8577
rect 1197 -8604 1215 -8586
rect 1269 -8595 1287 -8577
rect 1323 -8604 1341 -8586
<< psubstratepcontact >>
rect 135 -1503 171 -1467
rect 135 -1593 171 -1557
rect 945 -1503 981 -1467
rect 945 -1593 981 -1557
rect 1827 -1503 1863 -1467
rect 1827 -1593 1863 -1557
rect 135 -3600 171 -3564
rect 135 -3690 171 -3654
rect 945 -3600 981 -3564
rect 945 -3690 981 -3654
rect 1827 -3600 1863 -3564
rect 1827 -3690 1863 -3654
rect 135 -5715 171 -5679
rect 135 -5805 171 -5769
rect 945 -5715 981 -5679
rect 945 -5805 981 -5769
rect 1827 -5715 1863 -5679
rect 1827 -5805 1863 -5769
rect 135 -7650 171 -7614
rect 135 -7740 171 -7704
rect 945 -7650 981 -7614
rect 945 -7740 981 -7704
rect 1827 -7650 1863 -7614
rect 1827 -7740 1863 -7704
<< nsubstratencontact >>
rect 630 -1503 666 -1467
rect 630 -1593 666 -1557
rect 1440 -1503 1476 -1467
rect 1440 -1593 1476 -1557
rect 2322 -1503 2358 -1467
rect 2322 -1593 2358 -1557
rect 630 -3600 666 -3564
rect 630 -3690 666 -3654
rect 1440 -3600 1476 -3564
rect 1440 -3690 1476 -3654
rect 2322 -3600 2358 -3564
rect 2322 -3690 2358 -3654
rect 630 -5715 666 -5679
rect 630 -5805 666 -5769
rect 1440 -5715 1476 -5679
rect 1440 -5805 1476 -5769
rect 2322 -5715 2358 -5679
rect 2322 -5805 2358 -5769
rect 630 -7650 666 -7614
rect 630 -7740 666 -7704
rect 1440 -7650 1476 -7614
rect 1440 -7740 1476 -7704
rect 2322 -7650 2358 -7614
rect 2322 -7740 2358 -7704
<< polysilicon >>
rect 198 -1026 639 -1008
rect 198 -1116 216 -1026
rect 45 -1134 252 -1116
rect 306 -1134 315 -1116
rect 333 -1134 504 -1116
rect 567 -1134 594 -1116
rect -117 -3600 -99 -1521
rect 45 -1773 63 -1134
rect 333 -1287 351 -1134
rect 621 -1287 639 -1026
rect 1008 -1026 1449 -1008
rect 1008 -1116 1026 -1026
rect 855 -1134 1062 -1116
rect 1116 -1134 1125 -1116
rect 1143 -1134 1314 -1116
rect 1377 -1134 1404 -1116
rect 684 -1233 783 -1215
rect 90 -1305 252 -1287
rect 306 -1305 351 -1287
rect 468 -1305 504 -1287
rect 567 -1305 639 -1287
rect 90 -1647 108 -1305
rect 378 -1485 414 -1458
rect 189 -1503 252 -1485
rect 306 -1503 504 -1485
rect 567 -1503 612 -1485
rect 765 -1494 783 -1233
rect 387 -1566 405 -1503
rect 711 -1512 783 -1494
rect 216 -1575 405 -1566
rect 378 -1647 414 -1602
rect 90 -1665 252 -1647
rect 306 -1665 504 -1647
rect 567 -1665 612 -1647
rect 45 -1791 414 -1773
rect 711 -1791 729 -1512
rect 765 -1521 783 -1512
rect 783 -1539 792 -1521
rect 855 -1773 873 -1134
rect 1143 -1287 1161 -1134
rect 1431 -1287 1449 -1026
rect 1890 -1026 2331 -1008
rect 1890 -1116 1908 -1026
rect 1737 -1134 1944 -1116
rect 1998 -1134 2007 -1116
rect 2025 -1134 2196 -1116
rect 2259 -1134 2286 -1116
rect 1494 -1233 1620 -1215
rect 900 -1305 1062 -1287
rect 1116 -1305 1161 -1287
rect 1278 -1305 1314 -1287
rect 1377 -1305 1449 -1287
rect 900 -1647 918 -1305
rect 1188 -1485 1224 -1458
rect 999 -1503 1062 -1485
rect 1116 -1503 1314 -1485
rect 1377 -1503 1422 -1485
rect 1197 -1566 1215 -1503
rect 1602 -1521 1620 -1233
rect 1602 -1539 1647 -1521
rect 1044 -1575 1215 -1566
rect 1188 -1647 1224 -1602
rect 900 -1665 1062 -1647
rect 1116 -1665 1314 -1647
rect 1377 -1665 1422 -1647
rect 855 -1791 1224 -1773
rect 576 -1809 729 -1791
rect 576 -1917 594 -1809
rect 1251 -1872 1269 -1665
rect 1602 -1854 1620 -1539
rect 1665 -1539 1683 -1521
rect 1737 -1773 1755 -1134
rect 2025 -1287 2043 -1134
rect 2313 -1287 2331 -1026
rect 2376 -1242 2457 -1206
rect 1782 -1305 1944 -1287
rect 1998 -1305 2043 -1287
rect 2160 -1305 2196 -1287
rect 2259 -1305 2331 -1287
rect 1782 -1647 1800 -1305
rect 2070 -1485 2106 -1458
rect 1881 -1503 1944 -1485
rect 1998 -1503 2196 -1485
rect 2259 -1503 2304 -1485
rect 2079 -1566 2097 -1503
rect 1926 -1575 2097 -1566
rect 2070 -1611 2106 -1602
rect 2070 -1638 2079 -1611
rect 2097 -1638 2106 -1611
rect 2070 -1647 2106 -1638
rect 1782 -1665 1944 -1647
rect 1998 -1665 2196 -1647
rect 2259 -1665 2304 -1647
rect 1737 -1791 2106 -1773
rect 2133 -1809 2151 -1665
rect 2241 -1764 2556 -1746
rect 306 -1935 594 -1917
rect 684 -1890 1269 -1872
rect 1332 -1872 1620 -1854
rect 1710 -1827 2151 -1809
rect 306 -2169 324 -1935
rect 405 -2061 423 -2034
rect 567 -2061 585 -2034
rect 405 -2169 423 -2106
rect 306 -2187 423 -2169
rect 405 -2205 423 -2187
rect 567 -2178 585 -2106
rect 684 -2178 702 -1890
rect 864 -2025 882 -1908
rect 864 -2115 882 -2079
rect 873 -2142 882 -2115
rect 864 -2151 882 -2142
rect 567 -2196 702 -2178
rect 864 -2196 882 -2178
rect 567 -2205 585 -2196
rect 405 -2241 423 -2232
rect 567 -2241 585 -2232
rect 963 -2511 981 -2106
rect 1125 -2376 1143 -1971
rect 1206 -2214 1224 -1926
rect 1332 -2106 1350 -1872
rect 1431 -1998 1449 -1971
rect 1593 -1998 1611 -1971
rect 1431 -2106 1449 -2043
rect 1332 -2124 1449 -2106
rect 1431 -2142 1449 -2124
rect 1593 -2115 1611 -2043
rect 1710 -2115 1728 -1827
rect 1593 -2133 1728 -2115
rect 1593 -2142 1611 -2133
rect 1431 -2178 1449 -2169
rect 1593 -2178 1611 -2169
rect 1746 -2187 1764 -1854
rect 1890 -1962 1908 -1845
rect 1890 -2052 1908 -2016
rect 1899 -2079 1908 -2052
rect 1989 -2070 2025 -2043
rect 1890 -2088 1908 -2079
rect 1890 -2133 1908 -2115
rect 2007 -2259 2025 -2070
rect 1233 -2277 2025 -2259
rect 1080 -2421 1098 -2403
rect 1170 -2421 1188 -2403
rect 1080 -2511 1098 -2466
rect 963 -2529 1098 -2511
rect 1080 -2556 1098 -2529
rect 1170 -2538 1188 -2466
rect 1233 -2538 1251 -2277
rect 1296 -2421 1314 -2403
rect 1170 -2547 1251 -2538
rect 1296 -2511 1314 -2466
rect 1305 -2529 1314 -2511
rect 1170 -2556 1188 -2547
rect 1296 -2556 1314 -2529
rect 1080 -2592 1098 -2583
rect 1170 -2592 1188 -2583
rect 1296 -2592 1314 -2583
rect 2538 -3060 2556 -1764
rect 2538 -3087 2970 -3060
rect 198 -3123 639 -3105
rect 198 -3213 216 -3123
rect -117 -5715 -99 -3618
rect 45 -3231 252 -3213
rect 306 -3231 315 -3213
rect 333 -3231 504 -3213
rect 567 -3231 594 -3213
rect 45 -3870 63 -3231
rect 333 -3384 351 -3231
rect 621 -3384 639 -3123
rect 1008 -3123 1449 -3105
rect 1008 -3213 1026 -3123
rect 855 -3231 1062 -3213
rect 1116 -3231 1125 -3213
rect 1143 -3231 1314 -3213
rect 1377 -3231 1404 -3213
rect 684 -3330 783 -3312
rect 90 -3402 252 -3384
rect 306 -3402 351 -3384
rect 468 -3402 504 -3384
rect 567 -3402 639 -3384
rect 90 -3744 108 -3402
rect 378 -3582 414 -3555
rect 189 -3600 252 -3582
rect 306 -3600 504 -3582
rect 567 -3600 612 -3582
rect 765 -3591 783 -3330
rect 387 -3663 405 -3600
rect 711 -3609 783 -3591
rect 207 -3672 405 -3663
rect 378 -3744 414 -3699
rect 90 -3762 252 -3744
rect 306 -3762 504 -3744
rect 567 -3762 612 -3744
rect 45 -3888 414 -3870
rect 711 -3888 729 -3609
rect 765 -3618 783 -3609
rect 783 -3636 792 -3618
rect 855 -3870 873 -3231
rect 1143 -3384 1161 -3231
rect 1431 -3384 1449 -3123
rect 1890 -3123 2331 -3105
rect 1890 -3213 1908 -3123
rect 1737 -3231 1944 -3213
rect 1998 -3231 2007 -3213
rect 2025 -3231 2196 -3213
rect 2259 -3231 2286 -3213
rect 1494 -3330 1620 -3312
rect 900 -3402 1062 -3384
rect 1116 -3402 1161 -3384
rect 1278 -3402 1314 -3384
rect 1377 -3402 1449 -3384
rect 900 -3744 918 -3402
rect 1188 -3582 1224 -3555
rect 999 -3600 1062 -3582
rect 1116 -3600 1314 -3582
rect 1377 -3600 1422 -3582
rect 1197 -3663 1215 -3600
rect 1602 -3618 1620 -3330
rect 1602 -3636 1647 -3618
rect 1044 -3672 1215 -3663
rect 1188 -3744 1224 -3699
rect 900 -3762 1062 -3744
rect 1116 -3762 1314 -3744
rect 1377 -3762 1422 -3744
rect 855 -3888 1224 -3870
rect 576 -3906 729 -3888
rect 576 -4014 594 -3906
rect 1251 -3969 1269 -3762
rect 1602 -3951 1620 -3636
rect 1665 -3636 1683 -3618
rect 1737 -3870 1755 -3231
rect 2025 -3384 2043 -3231
rect 2313 -3384 2331 -3123
rect 2376 -3339 2457 -3303
rect 1782 -3402 1944 -3384
rect 1998 -3402 2043 -3384
rect 2160 -3402 2196 -3384
rect 2259 -3402 2331 -3384
rect 1782 -3744 1800 -3402
rect 2070 -3582 2106 -3555
rect 1881 -3600 1944 -3582
rect 1998 -3600 2196 -3582
rect 2259 -3600 2304 -3582
rect 2079 -3663 2097 -3600
rect 1926 -3672 2097 -3663
rect 2070 -3726 2079 -3699
rect 2097 -3726 2106 -3699
rect 2070 -3744 2106 -3726
rect 1782 -3762 1944 -3744
rect 1998 -3762 2196 -3744
rect 2259 -3762 2304 -3744
rect 1737 -3888 2106 -3870
rect 2133 -3906 2151 -3762
rect 2250 -3852 2826 -3834
rect 306 -4032 594 -4014
rect 684 -3987 1269 -3969
rect 1332 -3969 1620 -3951
rect 1710 -3924 2151 -3906
rect 306 -4266 324 -4032
rect 405 -4158 423 -4131
rect 567 -4158 585 -4131
rect 405 -4266 423 -4203
rect 306 -4284 423 -4266
rect 405 -4302 423 -4284
rect 567 -4275 585 -4203
rect 684 -4275 702 -3987
rect 864 -4122 882 -4005
rect 864 -4212 882 -4176
rect 873 -4239 882 -4212
rect 864 -4248 882 -4239
rect 567 -4293 702 -4275
rect 864 -4293 882 -4275
rect 567 -4302 585 -4293
rect 405 -4338 423 -4329
rect 567 -4338 585 -4329
rect 963 -4608 981 -4203
rect 1125 -4473 1143 -4068
rect 1206 -4311 1224 -4023
rect 1332 -4203 1350 -3969
rect 1431 -4095 1449 -4068
rect 1593 -4095 1611 -4068
rect 1431 -4203 1449 -4140
rect 1332 -4221 1449 -4203
rect 1431 -4239 1449 -4221
rect 1593 -4212 1611 -4140
rect 1710 -4212 1728 -3924
rect 1593 -4230 1728 -4212
rect 1593 -4239 1611 -4230
rect 1431 -4275 1449 -4266
rect 1593 -4275 1611 -4266
rect 1746 -4284 1764 -3951
rect 1890 -4059 1908 -3942
rect 1890 -4149 1908 -4113
rect 1899 -4176 1908 -4149
rect 1989 -4167 2025 -4140
rect 1890 -4185 1908 -4176
rect 1890 -4230 1908 -4212
rect 2007 -4356 2025 -4167
rect 1233 -4374 2025 -4356
rect 1080 -4518 1098 -4500
rect 1170 -4518 1188 -4500
rect 1080 -4608 1098 -4563
rect 963 -4626 1098 -4608
rect 1080 -4653 1098 -4626
rect 1170 -4635 1188 -4563
rect 1233 -4635 1251 -4374
rect 1296 -4518 1314 -4500
rect 1170 -4644 1251 -4635
rect 1296 -4608 1314 -4563
rect 1305 -4626 1314 -4608
rect 1170 -4653 1188 -4644
rect 1296 -4653 1314 -4626
rect 1080 -4689 1098 -4680
rect 1170 -4689 1188 -4680
rect 1296 -4689 1314 -4680
rect 198 -5238 639 -5220
rect 198 -5328 216 -5238
rect -117 -6570 -99 -5733
rect 45 -5346 252 -5328
rect 306 -5346 315 -5328
rect 333 -5346 504 -5328
rect 567 -5346 594 -5328
rect 45 -5985 63 -5346
rect 333 -5499 351 -5346
rect 621 -5499 639 -5238
rect 1008 -5238 1449 -5220
rect 1008 -5328 1026 -5238
rect 855 -5346 1062 -5328
rect 1116 -5346 1125 -5328
rect 1143 -5346 1314 -5328
rect 1377 -5346 1404 -5328
rect 684 -5445 783 -5427
rect 90 -5517 252 -5499
rect 306 -5517 351 -5499
rect 468 -5517 504 -5499
rect 567 -5517 639 -5499
rect 90 -5859 108 -5517
rect 378 -5697 414 -5670
rect 189 -5715 252 -5697
rect 306 -5715 504 -5697
rect 567 -5715 612 -5697
rect 765 -5706 783 -5445
rect 387 -5778 405 -5715
rect 711 -5724 783 -5706
rect 207 -5787 405 -5778
rect 378 -5859 414 -5814
rect 90 -5877 252 -5859
rect 306 -5877 504 -5859
rect 567 -5877 612 -5859
rect 45 -6003 414 -5985
rect 711 -6003 729 -5724
rect 765 -5733 783 -5724
rect 783 -5751 792 -5733
rect 855 -5985 873 -5346
rect 1143 -5499 1161 -5346
rect 1431 -5499 1449 -5238
rect 1890 -5238 2331 -5220
rect 1890 -5328 1908 -5238
rect 1737 -5346 1944 -5328
rect 1998 -5346 2007 -5328
rect 2025 -5346 2196 -5328
rect 2259 -5346 2286 -5328
rect 1494 -5445 1620 -5427
rect 900 -5517 1062 -5499
rect 1116 -5517 1161 -5499
rect 1278 -5517 1314 -5499
rect 1377 -5517 1449 -5499
rect 900 -5859 918 -5517
rect 1188 -5697 1224 -5670
rect 999 -5715 1062 -5697
rect 1116 -5715 1314 -5697
rect 1377 -5715 1422 -5697
rect 1197 -5778 1215 -5715
rect 1602 -5733 1620 -5445
rect 1602 -5751 1647 -5733
rect 1044 -5787 1215 -5778
rect 1188 -5859 1224 -5814
rect 900 -5877 1062 -5859
rect 1116 -5877 1314 -5859
rect 1377 -5877 1422 -5859
rect 855 -6003 1224 -5985
rect 576 -6021 729 -6003
rect 576 -6129 594 -6021
rect 1251 -6084 1269 -5877
rect 1602 -6066 1620 -5751
rect 1665 -5751 1683 -5733
rect 1737 -5985 1755 -5346
rect 2025 -5499 2043 -5346
rect 2313 -5499 2331 -5238
rect 2376 -5454 2457 -5418
rect 1782 -5517 1944 -5499
rect 1998 -5517 2043 -5499
rect 2160 -5517 2196 -5499
rect 2259 -5517 2331 -5499
rect 1782 -5859 1800 -5517
rect 2070 -5697 2106 -5670
rect 1881 -5715 1944 -5697
rect 1998 -5715 2196 -5697
rect 2259 -5715 2304 -5697
rect 2079 -5778 2097 -5715
rect 1926 -5787 2097 -5778
rect 2070 -5823 2106 -5814
rect 2070 -5841 2079 -5823
rect 2097 -5841 2106 -5823
rect 2070 -5859 2106 -5841
rect 1782 -5877 1944 -5859
rect 1998 -5877 2196 -5859
rect 2259 -5877 2304 -5859
rect 1737 -6003 2106 -5985
rect 2133 -6021 2151 -5877
rect 306 -6147 594 -6129
rect 684 -6102 1269 -6084
rect 1332 -6084 1620 -6066
rect 1710 -6039 2151 -6021
rect 306 -6381 324 -6147
rect 405 -6273 423 -6246
rect 567 -6273 585 -6246
rect 405 -6381 423 -6318
rect 306 -6399 423 -6381
rect 405 -6417 423 -6399
rect 567 -6390 585 -6318
rect 684 -6390 702 -6102
rect 864 -6237 882 -6120
rect 864 -6327 882 -6291
rect 873 -6354 882 -6327
rect 864 -6363 882 -6354
rect 567 -6408 702 -6390
rect 864 -6408 882 -6390
rect 567 -6417 585 -6408
rect 405 -6453 423 -6444
rect 567 -6453 585 -6444
rect -117 -6588 27 -6570
rect 9 -7578 27 -6588
rect 963 -6723 981 -6318
rect 1125 -6588 1143 -6183
rect 1206 -6426 1224 -6138
rect 1332 -6318 1350 -6084
rect 1431 -6210 1449 -6183
rect 1593 -6210 1611 -6183
rect 1431 -6318 1449 -6255
rect 1332 -6336 1449 -6318
rect 1431 -6354 1449 -6336
rect 1593 -6327 1611 -6255
rect 1710 -6327 1728 -6039
rect 1593 -6345 1728 -6327
rect 1593 -6354 1611 -6345
rect 1431 -6390 1449 -6381
rect 1593 -6390 1611 -6381
rect 1746 -6399 1764 -6066
rect 1890 -6174 1908 -6057
rect 1890 -6264 1908 -6228
rect 1899 -6291 1908 -6264
rect 1989 -6282 2025 -6255
rect 1890 -6300 1908 -6291
rect 1890 -6345 1908 -6327
rect 2007 -6471 2025 -6282
rect 1233 -6489 2025 -6471
rect 1080 -6633 1098 -6615
rect 1170 -6633 1188 -6615
rect 1080 -6723 1098 -6678
rect 963 -6741 1098 -6723
rect 1080 -6768 1098 -6741
rect 1170 -6750 1188 -6678
rect 1233 -6750 1251 -6489
rect 1296 -6633 1314 -6615
rect 1170 -6759 1251 -6750
rect 1296 -6723 1314 -6678
rect 2808 -6723 2826 -3852
rect 2952 -4608 2970 -3087
rect 1305 -6741 1314 -6723
rect 1368 -6741 2826 -6723
rect 1170 -6768 1188 -6759
rect 1296 -6768 1314 -6741
rect 1080 -6804 1098 -6795
rect 1170 -6804 1188 -6795
rect 1296 -6804 1314 -6795
rect 198 -7173 639 -7155
rect 198 -7263 216 -7173
rect 9 -7614 27 -7596
rect 45 -7281 252 -7263
rect 306 -7281 315 -7263
rect 333 -7281 504 -7263
rect 567 -7281 594 -7263
rect 45 -7920 63 -7281
rect 333 -7434 351 -7281
rect 621 -7434 639 -7173
rect 1008 -7173 1449 -7155
rect 1008 -7263 1026 -7173
rect 855 -7281 1062 -7263
rect 1116 -7281 1125 -7263
rect 1143 -7281 1314 -7263
rect 1377 -7281 1404 -7263
rect 684 -7380 783 -7362
rect 90 -7452 252 -7434
rect 306 -7452 351 -7434
rect 468 -7452 504 -7434
rect 567 -7452 639 -7434
rect 90 -7794 108 -7452
rect 378 -7632 414 -7605
rect 189 -7650 252 -7632
rect 306 -7650 504 -7632
rect 567 -7650 612 -7632
rect 765 -7641 783 -7380
rect 207 -7713 225 -7677
rect 387 -7713 405 -7650
rect 711 -7659 783 -7641
rect 207 -7722 405 -7713
rect 378 -7794 414 -7749
rect 90 -7812 252 -7794
rect 306 -7812 504 -7794
rect 567 -7812 612 -7794
rect 45 -7938 414 -7920
rect 711 -7938 729 -7659
rect 765 -7668 783 -7659
rect 783 -7686 792 -7668
rect 855 -7920 873 -7281
rect 1143 -7434 1161 -7281
rect 1431 -7434 1449 -7173
rect 1890 -7173 2331 -7155
rect 1890 -7263 1908 -7173
rect 1737 -7281 1944 -7263
rect 1998 -7281 2007 -7263
rect 2025 -7281 2196 -7263
rect 2259 -7281 2286 -7263
rect 1494 -7380 1620 -7362
rect 900 -7452 1062 -7434
rect 1116 -7452 1161 -7434
rect 1278 -7452 1314 -7434
rect 1377 -7452 1449 -7434
rect 900 -7794 918 -7452
rect 1188 -7632 1224 -7605
rect 999 -7650 1062 -7632
rect 1116 -7650 1314 -7632
rect 1377 -7650 1422 -7632
rect 1197 -7713 1215 -7650
rect 1602 -7668 1620 -7380
rect 1602 -7686 1647 -7668
rect 1044 -7722 1215 -7713
rect 1188 -7794 1224 -7749
rect 900 -7812 1062 -7794
rect 1116 -7812 1314 -7794
rect 1377 -7812 1422 -7794
rect 855 -7938 1224 -7920
rect 576 -7956 729 -7938
rect 576 -8064 594 -7956
rect 1251 -8019 1269 -7812
rect 1602 -8001 1620 -7686
rect 1665 -7686 1683 -7668
rect 1737 -7920 1755 -7281
rect 2025 -7434 2043 -7281
rect 2313 -7434 2331 -7173
rect 2376 -7389 2457 -7353
rect 1782 -7452 1944 -7434
rect 1998 -7452 2043 -7434
rect 2160 -7452 2196 -7434
rect 2259 -7452 2331 -7434
rect 1782 -7794 1800 -7452
rect 2070 -7632 2106 -7605
rect 1881 -7650 1944 -7632
rect 1998 -7650 2196 -7632
rect 2259 -7650 2304 -7632
rect 2079 -7713 2097 -7650
rect 1926 -7722 2097 -7713
rect 2070 -7758 2106 -7749
rect 2070 -7776 2079 -7758
rect 2097 -7776 2106 -7758
rect 2070 -7794 2106 -7776
rect 1782 -7812 1944 -7794
rect 1998 -7812 2196 -7794
rect 2259 -7812 2304 -7794
rect 1737 -7938 2106 -7920
rect 2133 -7956 2151 -7812
rect 306 -8082 594 -8064
rect 684 -8037 1269 -8019
rect 1332 -8019 1620 -8001
rect 1710 -7974 2151 -7956
rect 306 -8316 324 -8082
rect 405 -8208 423 -8181
rect 567 -8208 585 -8181
rect 405 -8316 423 -8253
rect 306 -8334 423 -8316
rect 405 -8352 423 -8334
rect 567 -8325 585 -8253
rect 684 -8325 702 -8037
rect 864 -8172 882 -8055
rect 864 -8262 882 -8226
rect 873 -8289 882 -8262
rect 864 -8298 882 -8289
rect 567 -8343 702 -8325
rect 864 -8343 882 -8325
rect 567 -8352 585 -8343
rect 405 -8388 423 -8379
rect 567 -8388 585 -8379
rect 963 -8658 981 -8253
rect 1125 -8523 1143 -8118
rect 1206 -8361 1224 -8073
rect 1332 -8253 1350 -8019
rect 1431 -8145 1449 -8118
rect 1593 -8145 1611 -8118
rect 1431 -8253 1449 -8190
rect 1332 -8271 1449 -8253
rect 1431 -8289 1449 -8271
rect 1593 -8262 1611 -8190
rect 1710 -8262 1728 -7974
rect 1593 -8280 1728 -8262
rect 1593 -8289 1611 -8280
rect 1431 -8325 1449 -8316
rect 1593 -8325 1611 -8316
rect 1746 -8334 1764 -8001
rect 1890 -8109 1908 -7992
rect 1890 -8199 1908 -8163
rect 1899 -8226 1908 -8199
rect 1989 -8217 2025 -8190
rect 1890 -8235 1908 -8226
rect 1890 -8280 1908 -8262
rect 2007 -8406 2025 -8217
rect 1233 -8424 2025 -8406
rect 1080 -8568 1098 -8550
rect 1170 -8568 1188 -8550
rect 1080 -8658 1098 -8613
rect 963 -8676 1098 -8658
rect 1080 -8703 1098 -8676
rect 1170 -8685 1188 -8613
rect 1233 -8685 1251 -8424
rect 1296 -8568 1314 -8550
rect 1170 -8694 1251 -8685
rect 1296 -8658 1314 -8613
rect 1305 -8676 1314 -8658
rect 1170 -8703 1188 -8694
rect 1296 -8703 1314 -8676
rect 1080 -8739 1098 -8730
rect 1170 -8739 1188 -8730
rect 1296 -8739 1314 -8730
<< polycontact >>
rect -117 -1521 -99 -1503
rect 648 -1233 684 -1215
rect 378 -1458 414 -1422
rect 198 -1575 216 -1548
rect 378 -1773 414 -1737
rect 765 -1539 783 -1521
rect 1458 -1233 1494 -1215
rect 1188 -1458 1224 -1422
rect 1017 -1584 1044 -1557
rect 1188 -1773 1224 -1737
rect 1647 -1548 1665 -1521
rect 2340 -1251 2376 -1206
rect 2070 -1458 2106 -1422
rect 1899 -1584 1926 -1557
rect 2079 -1638 2097 -1611
rect 2070 -1773 2106 -1737
rect 2214 -1764 2241 -1746
rect 1197 -1926 1224 -1908
rect 1125 -1971 1143 -1953
rect 846 -2142 873 -2115
rect 927 -2133 963 -2106
rect 1746 -1854 1764 -1836
rect 1872 -2079 1899 -2052
rect 1953 -2070 1989 -2043
rect 1746 -2205 1764 -2187
rect 1206 -2232 1224 -2214
rect 1125 -2394 1143 -2376
rect 1296 -2529 1305 -2511
rect -117 -3618 -99 -3600
rect 648 -3330 684 -3312
rect 378 -3555 414 -3519
rect 189 -3672 207 -3645
rect 378 -3870 414 -3834
rect 765 -3636 783 -3618
rect 1458 -3330 1494 -3312
rect 1188 -3555 1224 -3519
rect 1017 -3681 1044 -3654
rect 1188 -3870 1224 -3834
rect 1647 -3645 1665 -3618
rect 2340 -3348 2376 -3303
rect 2070 -3555 2106 -3519
rect 1899 -3681 1926 -3654
rect 2079 -3726 2097 -3699
rect 2070 -3870 2106 -3834
rect 2214 -3852 2250 -3834
rect 1197 -4023 1224 -4005
rect 1125 -4068 1143 -4050
rect 846 -4239 873 -4212
rect 927 -4230 963 -4203
rect 1746 -3951 1764 -3933
rect 1872 -4176 1899 -4149
rect 1953 -4167 1989 -4140
rect 1746 -4302 1764 -4284
rect 1206 -4329 1224 -4311
rect 1125 -4491 1143 -4473
rect 1296 -4626 1305 -4608
rect -117 -5733 -99 -5715
rect 648 -5445 684 -5427
rect 378 -5670 414 -5634
rect 189 -5787 207 -5760
rect 378 -5985 414 -5949
rect 765 -5751 783 -5733
rect 1458 -5445 1494 -5427
rect 1188 -5670 1224 -5634
rect 1017 -5796 1044 -5769
rect 1188 -5985 1224 -5949
rect 1647 -5760 1665 -5733
rect 2340 -5463 2376 -5418
rect 2070 -5670 2106 -5634
rect 1899 -5796 1926 -5769
rect 2079 -5841 2097 -5823
rect 2070 -5985 2106 -5949
rect 1197 -6138 1224 -6120
rect 1125 -6183 1143 -6165
rect 846 -6354 873 -6327
rect 927 -6345 963 -6318
rect 1746 -6066 1764 -6048
rect 1872 -6291 1899 -6264
rect 1953 -6282 1989 -6255
rect 1746 -6417 1764 -6399
rect 1206 -6444 1224 -6426
rect 1125 -6606 1143 -6588
rect 2943 -4626 2970 -4608
rect 1296 -6741 1305 -6723
rect 1332 -6741 1368 -6723
rect 9 -7596 27 -7578
rect 9 -7641 27 -7614
rect 648 -7380 684 -7362
rect 378 -7605 414 -7569
rect 207 -7677 225 -7659
rect 378 -7920 414 -7884
rect 765 -7686 783 -7668
rect 1458 -7380 1494 -7362
rect 1188 -7605 1224 -7569
rect 1017 -7731 1044 -7704
rect 1188 -7920 1224 -7884
rect 1647 -7695 1665 -7668
rect 2340 -7398 2376 -7353
rect 2070 -7605 2106 -7569
rect 1899 -7731 1926 -7704
rect 2079 -7776 2097 -7758
rect 2070 -7920 2106 -7884
rect 1197 -8073 1224 -8055
rect 1125 -8118 1143 -8100
rect 846 -8289 873 -8262
rect 927 -8280 963 -8253
rect 1746 -8001 1764 -7983
rect 1872 -8226 1899 -8199
rect 1953 -8217 1989 -8190
rect 1746 -8352 1764 -8334
rect 1206 -8379 1224 -8361
rect 1125 -8541 1143 -8523
rect 1296 -8676 1305 -8658
<< metal1 >>
rect 297 -1107 513 -1071
rect 549 -1107 729 -1071
rect 1107 -1107 1323 -1071
rect 1359 -1107 1539 -1071
rect 1989 -1107 2205 -1071
rect 2241 -1107 2421 -1071
rect 297 -1179 513 -1143
rect 549 -1179 684 -1143
rect 648 -1215 684 -1179
rect 135 -1278 261 -1242
rect 297 -1278 513 -1242
rect 135 -1377 171 -1278
rect 648 -1314 684 -1233
rect 297 -1350 513 -1314
rect 549 -1350 684 -1314
rect 693 -1377 729 -1107
rect 1107 -1179 1323 -1143
rect 1359 -1179 1494 -1143
rect 1458 -1215 1494 -1179
rect 135 -1413 360 -1377
rect 135 -1467 261 -1431
rect -99 -1521 -63 -1503
rect 135 -1530 171 -1503
rect -18 -1548 171 -1530
rect -18 -2250 0 -1548
rect 135 -1557 171 -1548
rect 324 -1512 360 -1413
rect 378 -1413 729 -1377
rect 945 -1278 1071 -1242
rect 1107 -1278 1323 -1242
rect 945 -1377 981 -1278
rect 1458 -1314 1494 -1233
rect 1107 -1350 1323 -1314
rect 1359 -1350 1494 -1314
rect 1503 -1377 1539 -1107
rect 1989 -1179 2205 -1143
rect 2241 -1179 2376 -1143
rect 2340 -1206 2376 -1179
rect 945 -1413 1170 -1377
rect 378 -1422 414 -1413
rect 549 -1467 666 -1431
rect 198 -1548 216 -1530
rect 297 -1548 513 -1512
rect 630 -1530 666 -1503
rect 945 -1467 1071 -1431
rect 630 -1548 756 -1530
rect 783 -1539 837 -1521
rect 630 -1557 666 -1548
rect 135 -1629 261 -1593
rect 549 -1629 666 -1593
rect 297 -1710 513 -1674
rect 378 -1737 414 -1710
rect 738 -1998 756 -1548
rect 945 -1557 981 -1503
rect 1134 -1512 1170 -1413
rect 1188 -1413 1539 -1377
rect 1827 -1278 1953 -1242
rect 1989 -1278 2205 -1242
rect 1827 -1377 1863 -1278
rect 2340 -1314 2376 -1251
rect 1989 -1350 2205 -1314
rect 2241 -1350 2376 -1314
rect 2385 -1377 2421 -1107
rect 1827 -1413 2052 -1377
rect 1188 -1422 1224 -1413
rect 1359 -1467 1476 -1431
rect 1107 -1548 1323 -1512
rect 1440 -1521 1476 -1503
rect 1827 -1467 1953 -1431
rect 1827 -1521 1863 -1503
rect 2016 -1512 2052 -1413
rect 2070 -1413 2421 -1377
rect 2070 -1422 2106 -1413
rect 2241 -1467 2358 -1431
rect 1440 -1539 1557 -1521
rect 1017 -1557 1035 -1548
rect 1440 -1557 1476 -1539
rect 945 -1629 1071 -1593
rect 1359 -1629 1476 -1593
rect 1017 -1908 1035 -1629
rect 1107 -1710 1323 -1674
rect 1188 -1737 1224 -1710
rect 1017 -1926 1197 -1908
rect 1539 -1935 1557 -1539
rect 1665 -1548 1692 -1521
rect 1818 -1539 1863 -1521
rect 1827 -1557 1863 -1539
rect 1989 -1548 2205 -1512
rect 2322 -1521 2358 -1503
rect 2322 -1539 2349 -1521
rect 1899 -1557 1926 -1548
rect 2322 -1557 2358 -1539
rect 1827 -1629 1953 -1593
rect 1854 -1836 1872 -1629
rect 2241 -1629 2358 -1593
rect 1989 -1710 2205 -1674
rect 2070 -1737 2106 -1710
rect 2205 -1764 2214 -1746
rect 1764 -1854 1872 -1836
rect 2385 -1890 2403 -1539
rect 1854 -1908 2403 -1890
rect 1854 -1935 1881 -1908
rect 1404 -1953 1881 -1935
rect 828 -1971 1125 -1953
rect 1143 -1971 1422 -1953
rect 828 -1998 855 -1971
rect 378 -2016 855 -1998
rect 378 -2070 396 -2016
rect 531 -2070 549 -2016
rect 828 -2025 855 -2016
rect 1404 -2007 1422 -1971
rect 1557 -2007 1575 -1953
rect 1854 -1962 1881 -1953
rect 432 -2151 450 -2097
rect 594 -2151 612 -2088
rect 756 -2142 846 -2115
rect 756 -2151 774 -2142
rect 432 -2169 774 -2151
rect 900 -2151 927 -2061
rect 1458 -2088 1476 -2034
rect 1620 -2088 1638 -2025
rect 1782 -2079 1872 -2052
rect 1782 -2088 1800 -2079
rect 1458 -2106 1800 -2088
rect 1926 -2088 1953 -1998
rect 1620 -2142 1638 -2106
rect 594 -2205 612 -2169
rect 1854 -2151 1881 -2124
rect 828 -2214 855 -2187
rect 1404 -2187 1422 -2169
rect 1854 -2169 1953 -2151
rect 1854 -2187 1890 -2169
rect 1404 -2205 1746 -2187
rect 1764 -2205 1890 -2187
rect 1404 -2214 1422 -2205
rect 378 -2250 396 -2232
rect 828 -2232 1206 -2214
rect 1224 -2232 1422 -2214
rect 828 -2250 864 -2232
rect -369 -2268 864 -2250
rect -369 -4347 -351 -2268
rect 846 -2601 864 -2268
rect 1044 -2394 1125 -2376
rect 1143 -2394 1314 -2376
rect 1044 -2430 1062 -2394
rect 1269 -2430 1287 -2394
rect 1197 -2511 1215 -2457
rect 1323 -2511 1341 -2457
rect 1107 -2529 1296 -2511
rect 1323 -2529 1368 -2511
rect 1107 -2556 1125 -2529
rect 1197 -2556 1215 -2529
rect 1323 -2556 1341 -2529
rect 1053 -2601 1071 -2574
rect 1143 -2601 1161 -2574
rect 1269 -2601 1287 -2574
rect 846 -2619 1287 -2601
rect 297 -3204 513 -3168
rect 549 -3204 729 -3168
rect 1107 -3204 1323 -3168
rect 1359 -3204 1539 -3168
rect 1989 -3204 2205 -3168
rect 2241 -3204 2421 -3168
rect 297 -3276 513 -3240
rect 549 -3276 684 -3240
rect 648 -3312 684 -3276
rect 135 -3375 261 -3339
rect 297 -3375 513 -3339
rect 135 -3474 171 -3375
rect 648 -3411 684 -3330
rect 297 -3447 513 -3411
rect 549 -3447 684 -3411
rect 693 -3474 729 -3204
rect 1107 -3276 1323 -3240
rect 1359 -3276 1494 -3240
rect 1458 -3312 1494 -3276
rect 135 -3510 360 -3474
rect 135 -3564 261 -3528
rect -99 -3618 -81 -3600
rect 135 -3627 171 -3600
rect 324 -3609 360 -3510
rect 378 -3510 729 -3474
rect 945 -3375 1071 -3339
rect 1107 -3375 1323 -3339
rect 945 -3474 981 -3375
rect 1458 -3411 1494 -3330
rect 1107 -3447 1323 -3411
rect 1359 -3447 1494 -3411
rect 1503 -3474 1539 -3204
rect 1989 -3276 2205 -3240
rect 2241 -3276 2376 -3240
rect 2340 -3303 2376 -3276
rect 945 -3510 1170 -3474
rect 378 -3519 414 -3510
rect 549 -3564 666 -3528
rect -18 -3645 171 -3627
rect -18 -4347 0 -3645
rect 135 -3654 171 -3645
rect 189 -3645 207 -3618
rect 297 -3645 513 -3609
rect 630 -3627 666 -3600
rect 945 -3564 1071 -3528
rect 630 -3645 756 -3627
rect 783 -3636 837 -3618
rect 630 -3654 666 -3645
rect 135 -3726 261 -3690
rect 549 -3726 666 -3690
rect 297 -3807 513 -3771
rect 378 -3834 414 -3807
rect 738 -4095 756 -3645
rect 945 -3654 981 -3600
rect 1134 -3609 1170 -3510
rect 1188 -3510 1539 -3474
rect 1827 -3375 1953 -3339
rect 1989 -3375 2205 -3339
rect 1827 -3474 1863 -3375
rect 2340 -3411 2376 -3348
rect 1989 -3447 2205 -3411
rect 2241 -3447 2376 -3411
rect 2385 -3474 2421 -3204
rect 1827 -3510 2052 -3474
rect 1188 -3519 1224 -3510
rect 1359 -3564 1476 -3528
rect 1107 -3645 1323 -3609
rect 1440 -3618 1476 -3600
rect 1827 -3564 1953 -3528
rect 1827 -3618 1863 -3600
rect 2016 -3609 2052 -3510
rect 2070 -3510 2421 -3474
rect 2070 -3519 2106 -3510
rect 2241 -3564 2358 -3528
rect 1440 -3636 1557 -3618
rect 1017 -3654 1035 -3645
rect 1440 -3654 1476 -3636
rect 945 -3726 1071 -3690
rect 1359 -3726 1476 -3690
rect 1017 -4005 1035 -3726
rect 1107 -3807 1323 -3771
rect 1188 -3834 1224 -3807
rect 1017 -4023 1197 -4005
rect 1539 -4032 1557 -3636
rect 1665 -3645 1692 -3618
rect 1818 -3636 1863 -3618
rect 1827 -3654 1863 -3636
rect 1989 -3645 2205 -3609
rect 2322 -3618 2358 -3600
rect 2322 -3636 2349 -3618
rect 2394 -3636 2403 -3618
rect 1899 -3654 1926 -3645
rect 2322 -3654 2358 -3636
rect 1827 -3726 1953 -3690
rect 2241 -3726 2358 -3690
rect 1854 -3933 1872 -3726
rect 2079 -3735 2097 -3726
rect 1989 -3807 2205 -3771
rect 2070 -3834 2106 -3807
rect 2196 -3852 2214 -3834
rect 1764 -3951 1872 -3933
rect 2385 -3987 2403 -3636
rect 1854 -4005 2403 -3987
rect 1854 -4032 1881 -4005
rect 1404 -4050 1881 -4032
rect 828 -4068 1125 -4050
rect 1143 -4068 1422 -4050
rect 828 -4095 855 -4068
rect 378 -4113 855 -4095
rect 378 -4167 396 -4113
rect 531 -4167 549 -4113
rect 828 -4122 855 -4113
rect 1404 -4104 1422 -4068
rect 1557 -4104 1575 -4050
rect 1854 -4059 1881 -4050
rect 432 -4248 450 -4194
rect 594 -4248 612 -4185
rect 756 -4239 846 -4212
rect 756 -4248 774 -4239
rect 432 -4266 774 -4248
rect 900 -4248 927 -4158
rect 1458 -4185 1476 -4131
rect 1620 -4185 1638 -4122
rect 1782 -4176 1872 -4149
rect 1782 -4185 1800 -4176
rect 1458 -4203 1800 -4185
rect 1926 -4185 1953 -4095
rect 1620 -4239 1638 -4203
rect 594 -4302 612 -4266
rect 1854 -4248 1881 -4221
rect 828 -4311 855 -4284
rect 1404 -4284 1422 -4266
rect 1854 -4266 1953 -4248
rect 1854 -4284 1890 -4266
rect 1404 -4302 1746 -4284
rect 1764 -4302 1890 -4284
rect 1404 -4311 1422 -4302
rect 378 -4347 396 -4329
rect 828 -4329 1206 -4311
rect 1224 -4329 1422 -4311
rect 828 -4347 864 -4329
rect -369 -4365 864 -4347
rect -369 -6462 -351 -4365
rect 846 -4698 864 -4365
rect 1044 -4491 1125 -4473
rect 1143 -4491 1314 -4473
rect 1044 -4527 1062 -4491
rect 1269 -4527 1287 -4491
rect 1197 -4608 1215 -4554
rect 1323 -4608 1341 -4554
rect 1107 -4626 1296 -4608
rect 1323 -4626 2943 -4608
rect 1107 -4653 1125 -4626
rect 1197 -4653 1215 -4626
rect 1323 -4653 1341 -4626
rect 1053 -4698 1071 -4671
rect 1143 -4698 1161 -4671
rect 1269 -4698 1287 -4671
rect 846 -4716 1287 -4698
rect 297 -5319 513 -5283
rect 549 -5319 729 -5283
rect 1107 -5319 1323 -5283
rect 1359 -5319 1539 -5283
rect 1989 -5319 2205 -5283
rect 2241 -5319 2421 -5283
rect 297 -5391 513 -5355
rect 549 -5391 684 -5355
rect 648 -5427 684 -5391
rect 135 -5490 261 -5454
rect 297 -5490 513 -5454
rect 135 -5589 171 -5490
rect 648 -5526 684 -5445
rect 297 -5562 513 -5526
rect 549 -5562 684 -5526
rect 693 -5589 729 -5319
rect 1107 -5391 1323 -5355
rect 1359 -5391 1494 -5355
rect 1458 -5427 1494 -5391
rect 135 -5625 360 -5589
rect 135 -5679 261 -5643
rect -99 -5733 -81 -5715
rect 135 -5742 171 -5715
rect 324 -5724 360 -5625
rect 378 -5625 729 -5589
rect 945 -5490 1071 -5454
rect 1107 -5490 1323 -5454
rect 945 -5589 981 -5490
rect 1458 -5526 1494 -5445
rect 1107 -5562 1323 -5526
rect 1359 -5562 1494 -5526
rect 1503 -5589 1539 -5319
rect 1989 -5391 2205 -5355
rect 2241 -5391 2376 -5355
rect 2340 -5418 2376 -5391
rect 945 -5625 1170 -5589
rect 378 -5634 414 -5625
rect 549 -5679 666 -5643
rect -18 -5760 171 -5742
rect -18 -6462 0 -5760
rect 135 -5769 171 -5760
rect 189 -5760 207 -5733
rect 297 -5760 513 -5724
rect 630 -5742 666 -5715
rect 945 -5679 1071 -5643
rect 630 -5760 756 -5742
rect 783 -5751 837 -5733
rect 630 -5769 666 -5760
rect 135 -5841 261 -5805
rect 549 -5841 666 -5805
rect 297 -5922 513 -5886
rect 378 -5949 414 -5922
rect 738 -6210 756 -5760
rect 945 -5769 981 -5715
rect 1134 -5724 1170 -5625
rect 1188 -5625 1539 -5589
rect 1827 -5490 1953 -5454
rect 1989 -5490 2205 -5454
rect 1827 -5589 1863 -5490
rect 2340 -5526 2376 -5463
rect 1989 -5562 2205 -5526
rect 2241 -5562 2376 -5526
rect 2385 -5589 2421 -5319
rect 1827 -5625 2052 -5589
rect 1188 -5634 1224 -5625
rect 1359 -5679 1476 -5643
rect 1107 -5760 1323 -5724
rect 1440 -5733 1476 -5715
rect 1827 -5679 1953 -5643
rect 1827 -5733 1863 -5715
rect 2016 -5724 2052 -5625
rect 2070 -5625 2421 -5589
rect 2070 -5634 2106 -5625
rect 2241 -5679 2358 -5643
rect 1440 -5751 1557 -5733
rect 1017 -5769 1035 -5760
rect 1440 -5769 1476 -5751
rect 945 -5841 1071 -5805
rect 1359 -5841 1476 -5805
rect 1017 -6120 1035 -5841
rect 1107 -5922 1323 -5886
rect 1188 -5949 1224 -5922
rect 1017 -6138 1197 -6120
rect 1539 -6147 1557 -5751
rect 1665 -5760 1692 -5733
rect 1818 -5751 1863 -5733
rect 1827 -5769 1863 -5751
rect 1989 -5760 2205 -5724
rect 2322 -5733 2358 -5715
rect 2322 -5751 2367 -5733
rect 1899 -5769 1926 -5760
rect 2322 -5769 2358 -5751
rect 1827 -5841 1953 -5805
rect 2241 -5841 2358 -5805
rect 1854 -6048 1872 -5841
rect 1989 -5922 2205 -5886
rect 2070 -5949 2106 -5922
rect 1764 -6066 1872 -6048
rect 2385 -6102 2403 -5751
rect 1854 -6120 2403 -6102
rect 1854 -6147 1881 -6120
rect 1404 -6165 1881 -6147
rect 828 -6183 1125 -6165
rect 1143 -6183 1422 -6165
rect 828 -6210 855 -6183
rect 378 -6228 855 -6210
rect 378 -6282 396 -6228
rect 531 -6282 549 -6228
rect 828 -6237 855 -6228
rect 1404 -6219 1422 -6183
rect 1557 -6219 1575 -6165
rect 1854 -6174 1881 -6165
rect 432 -6363 450 -6309
rect 594 -6363 612 -6300
rect 756 -6354 846 -6327
rect 756 -6363 774 -6354
rect 432 -6381 774 -6363
rect 900 -6363 927 -6273
rect 1458 -6300 1476 -6246
rect 1620 -6300 1638 -6237
rect 1782 -6291 1872 -6264
rect 1782 -6300 1800 -6291
rect 1458 -6318 1800 -6300
rect 1926 -6300 1953 -6210
rect 1620 -6354 1638 -6318
rect 594 -6417 612 -6381
rect 1854 -6363 1881 -6336
rect 828 -6426 855 -6399
rect 1404 -6399 1422 -6381
rect 1854 -6381 1953 -6363
rect 1854 -6399 1890 -6381
rect 1404 -6417 1746 -6399
rect 1764 -6417 1890 -6399
rect 1404 -6426 1422 -6417
rect 378 -6462 396 -6444
rect 828 -6444 1206 -6426
rect 1224 -6444 1422 -6426
rect 828 -6462 864 -6444
rect -369 -6480 864 -6462
rect -369 -8397 -351 -6480
rect 846 -6813 864 -6480
rect 1044 -6606 1125 -6588
rect 1143 -6606 1314 -6588
rect 1044 -6642 1062 -6606
rect 1269 -6642 1287 -6606
rect 1197 -6723 1215 -6669
rect 1323 -6723 1341 -6669
rect 1107 -6741 1296 -6723
rect 1323 -6741 1332 -6723
rect 1107 -6768 1125 -6741
rect 1197 -6768 1215 -6741
rect 1323 -6768 1341 -6741
rect 1053 -6813 1071 -6786
rect 1143 -6813 1161 -6786
rect 1269 -6813 1287 -6786
rect 846 -6831 1287 -6813
rect 297 -7254 513 -7218
rect 549 -7254 729 -7218
rect 1107 -7254 1323 -7218
rect 1359 -7254 1539 -7218
rect 1989 -7254 2205 -7218
rect 2241 -7254 2421 -7218
rect 297 -7326 513 -7290
rect 549 -7326 684 -7290
rect 648 -7362 684 -7326
rect 135 -7425 261 -7389
rect 297 -7425 513 -7389
rect 135 -7524 171 -7425
rect 648 -7461 684 -7380
rect 297 -7497 513 -7461
rect 549 -7497 684 -7461
rect 693 -7524 729 -7254
rect 1107 -7326 1323 -7290
rect 1359 -7326 1494 -7290
rect 1458 -7362 1494 -7326
rect 135 -7560 360 -7524
rect -45 -7596 9 -7578
rect 135 -7614 261 -7578
rect 9 -7659 27 -7641
rect 135 -7677 171 -7650
rect 324 -7659 360 -7560
rect 378 -7560 729 -7524
rect 945 -7425 1071 -7389
rect 1107 -7425 1323 -7389
rect 945 -7524 981 -7425
rect 1458 -7461 1494 -7380
rect 1107 -7497 1323 -7461
rect 1359 -7497 1494 -7461
rect 1503 -7524 1539 -7254
rect 1989 -7326 2205 -7290
rect 2241 -7326 2376 -7290
rect 2340 -7353 2376 -7326
rect 945 -7560 1170 -7524
rect 378 -7569 414 -7560
rect 549 -7614 666 -7578
rect 198 -7677 207 -7659
rect -18 -7695 171 -7677
rect 297 -7695 513 -7659
rect 630 -7677 666 -7650
rect 945 -7614 1071 -7578
rect 630 -7695 756 -7677
rect 783 -7686 837 -7668
rect -18 -8397 0 -7695
rect 135 -7704 171 -7695
rect 630 -7704 666 -7695
rect 135 -7776 261 -7740
rect 549 -7776 666 -7740
rect 297 -7857 513 -7821
rect 378 -7884 414 -7857
rect 738 -8145 756 -7695
rect 945 -7704 981 -7650
rect 1134 -7659 1170 -7560
rect 1188 -7560 1539 -7524
rect 1827 -7425 1953 -7389
rect 1989 -7425 2205 -7389
rect 1827 -7524 1863 -7425
rect 2340 -7461 2376 -7398
rect 1989 -7497 2205 -7461
rect 2241 -7497 2376 -7461
rect 2385 -7524 2421 -7254
rect 1827 -7560 2052 -7524
rect 1188 -7569 1224 -7560
rect 1359 -7614 1476 -7578
rect 1107 -7695 1323 -7659
rect 1440 -7668 1476 -7650
rect 1827 -7614 1953 -7578
rect 1827 -7668 1863 -7650
rect 2016 -7659 2052 -7560
rect 2070 -7560 2421 -7524
rect 2070 -7569 2106 -7560
rect 2241 -7614 2358 -7578
rect 1440 -7686 1557 -7668
rect 1017 -7704 1035 -7695
rect 1440 -7704 1476 -7686
rect 945 -7776 1071 -7740
rect 1359 -7776 1476 -7740
rect 1017 -8055 1035 -7776
rect 1107 -7857 1323 -7821
rect 1188 -7884 1224 -7857
rect 1017 -8073 1197 -8055
rect 1539 -8082 1557 -7686
rect 1665 -7695 1692 -7668
rect 1818 -7686 1863 -7668
rect 1827 -7704 1863 -7686
rect 1989 -7695 2205 -7659
rect 2322 -7668 2358 -7650
rect 2322 -7686 2367 -7668
rect 1899 -7704 1926 -7695
rect 2322 -7704 2358 -7686
rect 1827 -7776 1953 -7740
rect 2241 -7776 2358 -7740
rect 1854 -7983 1872 -7776
rect 1989 -7857 2205 -7821
rect 2070 -7884 2106 -7857
rect 1764 -8001 1872 -7983
rect 2385 -8037 2403 -7686
rect 1854 -8055 2403 -8037
rect 1854 -8082 1881 -8055
rect 1404 -8100 1881 -8082
rect 828 -8118 1125 -8100
rect 1143 -8118 1422 -8100
rect 828 -8145 855 -8118
rect 378 -8163 855 -8145
rect 378 -8217 396 -8163
rect 531 -8217 549 -8163
rect 828 -8172 855 -8163
rect 1404 -8154 1422 -8118
rect 1557 -8154 1575 -8100
rect 1854 -8109 1881 -8100
rect 432 -8298 450 -8244
rect 594 -8298 612 -8235
rect 756 -8289 846 -8262
rect 756 -8298 774 -8289
rect 432 -8316 774 -8298
rect 900 -8298 927 -8208
rect 1458 -8235 1476 -8181
rect 1620 -8235 1638 -8172
rect 1782 -8226 1872 -8199
rect 1782 -8235 1800 -8226
rect 1458 -8253 1800 -8235
rect 1926 -8235 1953 -8145
rect 1620 -8289 1638 -8253
rect 594 -8352 612 -8316
rect 1854 -8298 1881 -8271
rect 828 -8361 855 -8334
rect 1404 -8334 1422 -8316
rect 1854 -8316 1953 -8298
rect 1854 -8334 1890 -8316
rect 1404 -8352 1746 -8334
rect 1764 -8352 1890 -8334
rect 1404 -8361 1422 -8352
rect 378 -8397 396 -8379
rect 828 -8379 1206 -8361
rect 1224 -8379 1422 -8361
rect 828 -8397 864 -8379
rect -369 -8415 864 -8397
rect 846 -8748 864 -8415
rect 1044 -8541 1125 -8523
rect 1143 -8541 1314 -8523
rect 1044 -8577 1062 -8541
rect 1269 -8577 1287 -8541
rect 1197 -8658 1215 -8604
rect 1323 -8658 1341 -8604
rect 2745 -8658 2763 -5967
rect 1107 -8676 1296 -8658
rect 1323 -8676 2763 -8658
rect 1107 -8703 1125 -8676
rect 1197 -8703 1215 -8676
rect 1323 -8703 1341 -8676
rect 1053 -8748 1071 -8721
rect 1143 -8748 1161 -8721
rect 1269 -8748 1287 -8721
rect 846 -8766 1287 -8748
<< m2contact >>
rect -63 -1521 -27 -1503
rect 198 -1530 216 -1503
rect 837 -1539 864 -1512
rect 1017 -1548 1044 -1512
rect 1692 -1557 1728 -1521
rect 1899 -1548 1935 -1521
rect 2349 -1539 2403 -1521
rect 2079 -1665 2097 -1638
rect 2169 -1764 2205 -1746
rect -81 -3618 -45 -3600
rect 180 -3618 207 -3600
rect 837 -3636 864 -3609
rect 1017 -3645 1044 -3609
rect 1692 -3654 1728 -3618
rect 1899 -3645 1935 -3618
rect 2349 -3636 2394 -3618
rect 2079 -3762 2097 -3735
rect 2169 -3852 2196 -3834
rect -81 -5733 -54 -5715
rect 180 -5733 207 -5715
rect 837 -5751 864 -5724
rect 1017 -5760 1044 -5724
rect 1692 -5769 1728 -5733
rect 1899 -5760 1935 -5733
rect 2367 -5751 2403 -5733
rect 2079 -5868 2097 -5841
rect 2727 -5967 2763 -5949
rect -99 -7596 -45 -7578
rect 9 -7677 36 -7659
rect 180 -7677 198 -7659
rect 837 -7686 864 -7659
rect 1017 -7695 1044 -7659
rect 1692 -7704 1728 -7668
rect 1899 -7695 1935 -7668
rect 2367 -7686 2403 -7668
rect 2079 -7794 2097 -7776
<< metal2 >>
rect -27 -1521 198 -1503
rect 864 -1539 1017 -1521
rect 1728 -1548 1899 -1521
rect 2403 -1539 2871 -1521
rect 2079 -1638 2097 -1629
rect 2079 -1683 2097 -1665
rect 2079 -1701 2169 -1683
rect 2151 -1764 2169 -1701
rect -45 -3618 180 -3600
rect 864 -3636 1017 -3618
rect 2853 -3618 2871 -1539
rect 1728 -3645 1899 -3618
rect 2394 -3636 2871 -3618
rect 2079 -3780 2097 -3762
rect 2079 -3798 2169 -3780
rect 2151 -3852 2169 -3798
rect -54 -5733 180 -5715
rect 864 -5751 1017 -5733
rect 2853 -5733 2871 -3636
rect 1728 -5760 1899 -5733
rect 2403 -5751 2871 -5733
rect 2079 -5895 2097 -5868
rect 2079 -5913 2169 -5895
rect 2151 -5949 2169 -5913
rect 2151 -5967 2727 -5949
rect -180 -7596 -99 -7578
rect -180 -8793 -162 -7596
rect 36 -7677 180 -7659
rect 864 -7686 1017 -7668
rect 2853 -7668 2871 -5751
rect 1728 -7695 1899 -7668
rect 2403 -7686 2871 -7668
rect 2385 -7695 2403 -7686
rect 2079 -7830 2097 -7794
rect 2079 -7848 2169 -7830
rect 2151 -7911 2169 -7848
rect 2151 -7929 2475 -7911
rect 2457 -8793 2475 -7929
rect -180 -8811 2475 -8793
<< labels >>
rlabel polysilicon -108 -4221 -108 -4221 3 d1
rlabel polysilicon 396 -1629 396 -1629 1 b3_adsub
rlabel polysilicon 396 -3735 396 -3735 1 b2_adsub
rlabel polysilicon 396 -5841 396 -5841 1 b1_adsub
rlabel polysilicon 396 -7776 396 -7776 1 b0_adsub
rlabel polysilicon 1206 -1629 1206 -1629 1 a3_adsub
rlabel polysilicon 1206 -3726 1206 -3726 1 a2_adsub
rlabel polysilicon 1215 -5841 1215 -5841 1 a1_adsub
rlabel polysilicon 1206 -7776 1206 -7776 1 a0_adsub
rlabel polysilicon 2439 -7371 2439 -7371 7 sum0
rlabel metal1 1359 -8667 1359 -8667 1 carry0
rlabel polysilicon 2448 -5436 2448 -5436 1 sum1
rlabel polycontact 1350 -6732 1350 -6732 1 carry1
rlabel polysilicon 2430 -3321 2430 -3321 1 sum2
rlabel metal1 1350 -4617 1350 -4617 1 carry2
rlabel polysilicon 2439 -1224 2439 -1224 1 sum3
rlabel metal1 1350 -2520 1350 -2520 1 carry3
rlabel metal1 855 -8667 855 -8667 1 gnd
rlabel metal1 2142 -8046 2142 -8046 1 vdd
<< end >>
