magic
tech scmos
magscale 9 1
timestamp 1700920048
<< nwell >>
rect 46 83 67 89
rect -6 66 30 76
rect 46 71 63 83
rect 46 70 53 71
rect 55 70 63 71
rect 46 28 67 34
rect -6 11 30 21
rect 46 16 63 28
rect 46 15 53 16
rect 55 15 63 16
rect 46 -18 67 -12
rect -6 -35 30 -25
rect 46 -30 63 -18
rect 46 -31 53 -30
rect 55 -31 63 -30
rect 46 -77 67 -71
rect -6 -94 30 -84
rect 46 -89 63 -77
rect 46 -90 53 -89
rect 55 -90 63 -89
rect 46 -132 67 -126
rect -6 -149 30 -139
rect 46 -144 63 -132
rect 46 -145 53 -144
rect 55 -145 63 -144
rect 46 -187 67 -181
rect -6 -204 30 -194
rect 46 -199 63 -187
rect 46 -200 53 -199
rect 55 -200 63 -199
rect 46 -233 67 -227
rect -6 -250 30 -240
rect 46 -245 63 -233
rect 46 -246 53 -245
rect 55 -246 63 -245
rect 46 -292 67 -286
rect -6 -309 30 -299
rect 46 -304 63 -292
rect 46 -305 53 -304
rect 55 -305 63 -304
<< ntransistor >>
rect 53 61 55 64
rect 2 55 4 58
rect 20 55 22 58
rect 53 6 55 9
rect 2 0 4 3
rect 20 0 22 3
rect 53 -40 55 -37
rect 2 -46 4 -43
rect 20 -46 22 -43
rect 53 -99 55 -96
rect 2 -105 4 -102
rect 20 -105 22 -102
rect 53 -154 55 -151
rect 2 -160 4 -157
rect 20 -160 22 -157
rect 53 -209 55 -206
rect 2 -215 4 -212
rect 20 -215 22 -212
rect 53 -255 55 -252
rect 2 -261 4 -258
rect 20 -261 22 -258
rect 53 -314 55 -311
rect 2 -320 4 -317
rect 20 -320 22 -317
<< ptransistor >>
rect 2 69 4 74
rect 20 69 22 74
rect 53 72 55 78
rect 2 14 4 19
rect 20 14 22 19
rect 53 17 55 23
rect 2 -32 4 -27
rect 20 -32 22 -27
rect 53 -29 55 -23
rect 2 -91 4 -86
rect 20 -91 22 -86
rect 53 -88 55 -82
rect 2 -146 4 -141
rect 20 -146 22 -141
rect 53 -143 55 -137
rect 2 -201 4 -196
rect 20 -201 22 -196
rect 53 -198 55 -192
rect 2 -247 4 -242
rect 20 -247 22 -242
rect 53 -244 55 -238
rect 2 -306 4 -301
rect 20 -306 22 -301
rect 53 -303 55 -297
<< ndiffusion >>
rect 48 63 53 64
rect 48 61 49 63
rect 52 61 53 63
rect 55 61 57 64
rect 60 61 61 64
rect -2 57 2 58
rect -2 55 -1 57
rect 1 55 2 57
rect 4 55 20 58
rect 22 56 23 58
rect 25 56 26 58
rect 22 55 26 56
rect 48 8 53 9
rect 48 6 49 8
rect 52 6 53 8
rect 55 6 57 9
rect 60 6 61 9
rect -2 2 2 3
rect -2 0 -1 2
rect 1 0 2 2
rect 4 0 20 3
rect 22 1 23 3
rect 25 1 26 3
rect 22 0 26 1
rect 48 -38 53 -37
rect 48 -40 49 -38
rect 52 -40 53 -38
rect 55 -40 57 -37
rect 60 -40 61 -37
rect -2 -44 2 -43
rect -2 -46 -1 -44
rect 1 -46 2 -44
rect 4 -46 20 -43
rect 22 -45 23 -43
rect 25 -45 26 -43
rect 22 -46 26 -45
rect 48 -97 53 -96
rect 48 -99 49 -97
rect 52 -99 53 -97
rect 55 -99 57 -96
rect 60 -99 61 -96
rect -2 -103 2 -102
rect -2 -105 -1 -103
rect 1 -105 2 -103
rect 4 -105 20 -102
rect 22 -104 23 -102
rect 25 -104 26 -102
rect 22 -105 26 -104
rect 48 -152 53 -151
rect 48 -154 49 -152
rect 52 -154 53 -152
rect 55 -154 57 -151
rect 60 -154 61 -151
rect -2 -158 2 -157
rect -2 -160 -1 -158
rect 1 -160 2 -158
rect 4 -160 20 -157
rect 22 -159 23 -157
rect 25 -159 26 -157
rect 22 -160 26 -159
rect 48 -207 53 -206
rect 48 -209 49 -207
rect 52 -209 53 -207
rect 55 -209 57 -206
rect 60 -209 61 -206
rect -2 -213 2 -212
rect -2 -215 -1 -213
rect 1 -215 2 -213
rect 4 -215 20 -212
rect 22 -214 23 -212
rect 25 -214 26 -212
rect 22 -215 26 -214
rect 48 -253 53 -252
rect 48 -255 49 -253
rect 52 -255 53 -253
rect 55 -255 57 -252
rect 60 -255 61 -252
rect -2 -259 2 -258
rect -2 -261 -1 -259
rect 1 -261 2 -259
rect 4 -261 20 -258
rect 22 -260 23 -258
rect 25 -260 26 -258
rect 22 -261 26 -260
rect 48 -312 53 -311
rect 48 -314 49 -312
rect 52 -314 53 -312
rect 55 -314 57 -311
rect 60 -314 61 -311
rect -2 -318 2 -317
rect -2 -320 -1 -318
rect 1 -320 2 -318
rect 4 -320 20 -317
rect 22 -319 23 -317
rect 25 -319 26 -317
rect 22 -320 26 -319
<< pdiffusion >>
rect 48 75 49 78
rect 52 75 53 78
rect -2 73 2 74
rect -2 71 -1 73
rect 1 71 2 73
rect -2 69 2 71
rect 4 72 11 74
rect 4 70 5 72
rect 7 70 11 72
rect 4 69 11 70
rect 15 73 20 74
rect 15 71 16 73
rect 18 71 20 73
rect 15 69 20 71
rect 22 73 26 74
rect 22 71 23 73
rect 25 71 26 73
rect 48 72 53 75
rect 55 77 61 78
rect 55 74 57 77
rect 60 74 61 77
rect 55 72 61 74
rect 22 69 26 71
rect 48 20 49 23
rect 52 20 53 23
rect -2 18 2 19
rect -2 16 -1 18
rect 1 16 2 18
rect -2 14 2 16
rect 4 17 11 19
rect 4 15 5 17
rect 7 15 11 17
rect 4 14 11 15
rect 15 18 20 19
rect 15 16 16 18
rect 18 16 20 18
rect 15 14 20 16
rect 22 18 26 19
rect 22 16 23 18
rect 25 16 26 18
rect 48 17 53 20
rect 55 22 61 23
rect 55 19 57 22
rect 60 19 61 22
rect 55 17 61 19
rect 22 14 26 16
rect 48 -26 49 -23
rect 52 -26 53 -23
rect -2 -28 2 -27
rect -2 -30 -1 -28
rect 1 -30 2 -28
rect -2 -32 2 -30
rect 4 -29 11 -27
rect 4 -31 5 -29
rect 7 -31 11 -29
rect 4 -32 11 -31
rect 15 -28 20 -27
rect 15 -30 16 -28
rect 18 -30 20 -28
rect 15 -32 20 -30
rect 22 -28 26 -27
rect 22 -30 23 -28
rect 25 -30 26 -28
rect 48 -29 53 -26
rect 55 -24 61 -23
rect 55 -27 57 -24
rect 60 -27 61 -24
rect 55 -29 61 -27
rect 22 -32 26 -30
rect 48 -85 49 -82
rect 52 -85 53 -82
rect -2 -87 2 -86
rect -2 -89 -1 -87
rect 1 -89 2 -87
rect -2 -91 2 -89
rect 4 -88 11 -86
rect 4 -90 5 -88
rect 7 -90 11 -88
rect 4 -91 11 -90
rect 15 -87 20 -86
rect 15 -89 16 -87
rect 18 -89 20 -87
rect 15 -91 20 -89
rect 22 -87 26 -86
rect 22 -89 23 -87
rect 25 -89 26 -87
rect 48 -88 53 -85
rect 55 -83 61 -82
rect 55 -86 57 -83
rect 60 -86 61 -83
rect 55 -88 61 -86
rect 22 -91 26 -89
rect 48 -140 49 -137
rect 52 -140 53 -137
rect -2 -142 2 -141
rect -2 -144 -1 -142
rect 1 -144 2 -142
rect -2 -146 2 -144
rect 4 -143 11 -141
rect 4 -145 5 -143
rect 7 -145 11 -143
rect 4 -146 11 -145
rect 15 -142 20 -141
rect 15 -144 16 -142
rect 18 -144 20 -142
rect 15 -146 20 -144
rect 22 -142 26 -141
rect 22 -144 23 -142
rect 25 -144 26 -142
rect 48 -143 53 -140
rect 55 -138 61 -137
rect 55 -141 57 -138
rect 60 -141 61 -138
rect 55 -143 61 -141
rect 22 -146 26 -144
rect 48 -195 49 -192
rect 52 -195 53 -192
rect -2 -197 2 -196
rect -2 -199 -1 -197
rect 1 -199 2 -197
rect -2 -201 2 -199
rect 4 -198 11 -196
rect 4 -200 5 -198
rect 7 -200 11 -198
rect 4 -201 11 -200
rect 15 -197 20 -196
rect 15 -199 16 -197
rect 18 -199 20 -197
rect 15 -201 20 -199
rect 22 -197 26 -196
rect 22 -199 23 -197
rect 25 -199 26 -197
rect 48 -198 53 -195
rect 55 -193 61 -192
rect 55 -196 57 -193
rect 60 -196 61 -193
rect 55 -198 61 -196
rect 22 -201 26 -199
rect 48 -241 49 -238
rect 52 -241 53 -238
rect -2 -243 2 -242
rect -2 -245 -1 -243
rect 1 -245 2 -243
rect -2 -247 2 -245
rect 4 -244 11 -242
rect 4 -246 5 -244
rect 7 -246 11 -244
rect 4 -247 11 -246
rect 15 -243 20 -242
rect 15 -245 16 -243
rect 18 -245 20 -243
rect 15 -247 20 -245
rect 22 -243 26 -242
rect 22 -245 23 -243
rect 25 -245 26 -243
rect 48 -244 53 -241
rect 55 -239 61 -238
rect 55 -242 57 -239
rect 60 -242 61 -239
rect 55 -244 61 -242
rect 22 -247 26 -245
rect 48 -300 49 -297
rect 52 -300 53 -297
rect -2 -302 2 -301
rect -2 -304 -1 -302
rect 1 -304 2 -302
rect -2 -306 2 -304
rect 4 -303 11 -301
rect 4 -305 5 -303
rect 7 -305 11 -303
rect 4 -306 11 -305
rect 15 -302 20 -301
rect 15 -304 16 -302
rect 18 -304 20 -302
rect 15 -306 20 -304
rect 22 -302 26 -301
rect 22 -304 23 -302
rect 25 -304 26 -302
rect 48 -303 53 -300
rect 55 -298 61 -297
rect 55 -301 57 -298
rect 60 -301 61 -298
rect 55 -303 61 -301
rect 22 -306 26 -304
<< ndcontact >>
rect 49 60 52 63
rect 57 61 60 64
rect -1 55 1 57
rect 23 56 25 58
rect 49 5 52 8
rect 57 6 60 9
rect -1 0 1 2
rect 23 1 25 3
rect 49 -41 52 -38
rect 57 -40 60 -37
rect -1 -46 1 -44
rect 23 -45 25 -43
rect 49 -100 52 -97
rect 57 -99 60 -96
rect -1 -105 1 -103
rect 23 -104 25 -102
rect 49 -155 52 -152
rect 57 -154 60 -151
rect -1 -160 1 -158
rect 23 -159 25 -157
rect 49 -210 52 -207
rect 57 -209 60 -206
rect -1 -215 1 -213
rect 23 -214 25 -212
rect 49 -256 52 -253
rect 57 -255 60 -252
rect -1 -261 1 -259
rect 23 -260 25 -258
rect 49 -315 52 -312
rect 57 -314 60 -311
rect -1 -320 1 -318
rect 23 -319 25 -317
<< pdcontact >>
rect 49 75 52 78
rect -1 71 1 73
rect 5 70 7 72
rect 16 71 18 73
rect 23 71 25 73
rect 57 74 60 77
rect 49 20 52 23
rect -1 16 1 18
rect 5 15 7 17
rect 16 16 18 18
rect 23 16 25 18
rect 57 19 60 22
rect 49 -26 52 -23
rect -1 -30 1 -28
rect 5 -31 7 -29
rect 16 -30 18 -28
rect 23 -30 25 -28
rect 57 -27 60 -24
rect 49 -85 52 -82
rect -1 -89 1 -87
rect 5 -90 7 -88
rect 16 -89 18 -87
rect 23 -89 25 -87
rect 57 -86 60 -83
rect 49 -140 52 -137
rect -1 -144 1 -142
rect 5 -145 7 -143
rect 16 -144 18 -142
rect 23 -144 25 -142
rect 57 -141 60 -138
rect 49 -195 52 -192
rect -1 -199 1 -197
rect 5 -200 7 -198
rect 16 -199 18 -197
rect 23 -199 25 -197
rect 57 -196 60 -193
rect 49 -241 52 -238
rect -1 -245 1 -243
rect 5 -246 7 -244
rect 16 -245 18 -243
rect 23 -245 25 -243
rect 57 -242 60 -239
rect 49 -300 52 -297
rect -1 -304 1 -302
rect 5 -305 7 -303
rect 16 -304 18 -302
rect 23 -304 25 -302
rect 57 -301 60 -298
<< polysilicon >>
rect 53 78 55 91
rect 2 74 4 77
rect 20 74 22 77
rect 2 62 4 69
rect -17 60 4 62
rect -17 7 -15 60
rect 2 58 4 60
rect 20 58 22 69
rect 53 68 55 72
rect 54 65 55 68
rect 53 64 55 65
rect 53 59 55 61
rect 2 54 4 55
rect 20 54 22 55
rect 53 23 55 36
rect 2 19 4 22
rect 20 19 22 22
rect 2 7 4 14
rect -17 5 4 7
rect -17 -40 -15 5
rect 2 3 4 5
rect 20 3 22 14
rect 53 13 55 17
rect 54 10 55 13
rect 53 9 55 10
rect 53 4 55 6
rect 2 -1 4 0
rect 20 -1 22 0
rect 53 -23 55 -10
rect 2 -27 4 -24
rect 20 -27 22 -24
rect 2 -40 4 -32
rect -17 -42 4 -40
rect -17 -98 -15 -42
rect 2 -43 4 -42
rect 20 -43 22 -32
rect 53 -33 55 -29
rect 54 -36 55 -33
rect 53 -37 55 -36
rect 53 -42 55 -40
rect 2 -47 4 -46
rect 20 -47 22 -46
rect 53 -82 55 -69
rect 2 -86 4 -83
rect 20 -86 22 -83
rect 2 -98 4 -91
rect -17 -100 4 -98
rect -17 -153 -15 -100
rect 2 -102 4 -100
rect 20 -102 22 -91
rect 53 -92 55 -88
rect 54 -95 55 -92
rect 53 -96 55 -95
rect 53 -101 55 -99
rect 2 -106 4 -105
rect 20 -106 22 -105
rect 53 -137 55 -124
rect 2 -141 4 -138
rect 20 -141 22 -138
rect 2 -153 4 -146
rect -17 -155 4 -153
rect -17 -208 -15 -155
rect 2 -157 4 -155
rect 20 -157 22 -146
rect 53 -147 55 -143
rect 54 -150 55 -147
rect 53 -151 55 -150
rect 53 -156 55 -154
rect 2 -161 4 -160
rect 20 -161 22 -160
rect 53 -192 55 -179
rect 2 -196 4 -193
rect 20 -196 22 -193
rect 2 -208 4 -201
rect -17 -210 4 -208
rect -17 -255 -15 -210
rect 2 -212 4 -210
rect 20 -212 22 -201
rect 53 -202 55 -198
rect 54 -205 55 -202
rect 53 -206 55 -205
rect 53 -211 55 -209
rect 2 -216 4 -215
rect 20 -216 22 -215
rect 53 -238 55 -225
rect 2 -242 4 -239
rect 20 -242 22 -239
rect 2 -255 4 -247
rect -17 -257 4 -255
rect -17 -313 -15 -257
rect 2 -258 4 -257
rect 20 -258 22 -247
rect 53 -248 55 -244
rect 54 -251 55 -248
rect 53 -252 55 -251
rect 53 -257 55 -255
rect 2 -262 4 -261
rect 20 -262 22 -261
rect 53 -297 55 -284
rect 2 -301 4 -298
rect 20 -301 22 -298
rect 2 -313 4 -306
rect -17 -315 4 -313
rect 2 -317 4 -315
rect 20 -317 22 -306
rect 53 -307 55 -303
rect 54 -310 55 -307
rect 53 -311 55 -310
rect 53 -316 55 -314
rect 2 -321 4 -320
rect 20 -321 22 -320
<< polycontact >>
rect 51 65 54 68
rect 51 10 54 13
rect 51 -36 54 -33
rect 51 -95 54 -92
rect 51 -150 54 -147
rect 51 -205 54 -202
rect 51 -251 54 -248
rect 51 -310 54 -307
<< metal1 >>
rect 49 84 75 86
rect 49 81 52 84
rect -1 79 52 81
rect -1 73 1 79
rect 16 73 18 79
rect 49 78 52 79
rect 5 64 7 70
rect 23 64 25 71
rect 57 69 60 74
rect 41 65 51 68
rect 57 66 63 69
rect 41 64 43 65
rect 5 62 43 64
rect 57 64 60 66
rect 23 58 25 62
rect 49 57 52 60
rect -1 53 1 55
rect 49 55 60 57
rect 49 53 53 55
rect -13 51 53 53
rect -13 -2 -11 51
rect 73 31 75 84
rect 49 29 75 31
rect 49 26 52 29
rect -1 24 52 26
rect -1 18 1 24
rect 16 18 18 24
rect 49 23 52 24
rect 5 9 7 15
rect 23 9 25 16
rect 57 14 60 19
rect 41 10 51 13
rect 57 11 63 14
rect 41 9 43 10
rect 5 7 43 9
rect 57 9 60 11
rect 23 3 25 7
rect 49 2 52 5
rect -1 -2 1 0
rect 49 0 60 2
rect 49 -2 53 0
rect -13 -4 53 -2
rect -13 -48 -11 -4
rect 73 -15 75 29
rect 49 -17 75 -15
rect 49 -20 52 -17
rect -1 -22 52 -20
rect -1 -28 1 -22
rect 16 -28 18 -22
rect 49 -23 52 -22
rect 5 -37 7 -31
rect 23 -37 25 -30
rect 57 -32 60 -27
rect 41 -36 51 -33
rect 57 -35 63 -32
rect 41 -37 43 -36
rect 5 -39 43 -37
rect 57 -37 60 -35
rect 23 -43 25 -39
rect 49 -44 52 -41
rect -1 -48 1 -46
rect 49 -46 60 -44
rect 49 -48 53 -46
rect -13 -50 53 -48
rect -13 -107 -11 -50
rect 73 -74 75 -17
rect 49 -76 75 -74
rect 49 -79 52 -76
rect -1 -81 52 -79
rect -1 -87 1 -81
rect 16 -87 18 -81
rect 49 -82 52 -81
rect 5 -96 7 -90
rect 23 -96 25 -89
rect 57 -91 60 -86
rect 41 -95 51 -92
rect 57 -94 63 -91
rect 41 -96 43 -95
rect 5 -98 43 -96
rect 57 -96 60 -94
rect 23 -102 25 -98
rect 49 -103 52 -100
rect -1 -107 1 -105
rect 49 -105 60 -103
rect 49 -107 53 -105
rect -13 -109 53 -107
rect -13 -162 -11 -109
rect 73 -129 75 -76
rect 49 -131 75 -129
rect 49 -134 52 -131
rect -1 -136 52 -134
rect -1 -142 1 -136
rect 16 -142 18 -136
rect 49 -137 52 -136
rect 5 -151 7 -145
rect 23 -151 25 -144
rect 57 -146 60 -141
rect 41 -150 51 -147
rect 57 -149 63 -146
rect 41 -151 43 -150
rect 5 -153 43 -151
rect 57 -151 60 -149
rect 23 -157 25 -153
rect 49 -158 52 -155
rect -1 -162 1 -160
rect 49 -160 56 -158
rect 49 -162 53 -160
rect -13 -164 53 -162
rect -13 -217 -11 -164
rect 73 -184 75 -131
rect 49 -186 75 -184
rect 49 -189 52 -186
rect -1 -191 52 -189
rect -1 -197 1 -191
rect 16 -197 18 -191
rect 49 -192 52 -191
rect 5 -206 7 -200
rect 23 -206 25 -199
rect 57 -201 60 -196
rect 41 -205 51 -202
rect 57 -204 63 -201
rect 41 -206 43 -205
rect 5 -208 43 -206
rect 57 -206 60 -204
rect 23 -212 25 -208
rect 49 -213 52 -210
rect -1 -217 1 -215
rect 49 -215 60 -213
rect 49 -217 53 -215
rect -13 -219 53 -217
rect -13 -263 -11 -219
rect 73 -230 75 -186
rect 49 -232 75 -230
rect 49 -235 52 -232
rect -1 -237 52 -235
rect -1 -243 1 -237
rect 16 -243 18 -237
rect 49 -238 52 -237
rect 5 -252 7 -246
rect 23 -252 25 -245
rect 57 -247 60 -242
rect 41 -251 51 -248
rect 57 -250 63 -247
rect 41 -252 43 -251
rect 5 -254 43 -252
rect 57 -252 60 -250
rect 23 -258 25 -254
rect 49 -259 52 -256
rect -1 -263 1 -261
rect 49 -261 60 -259
rect 49 -263 53 -261
rect -13 -265 53 -263
rect -13 -322 -11 -265
rect 73 -289 75 -232
rect 49 -291 75 -289
rect 49 -294 52 -291
rect -1 -296 52 -294
rect -1 -302 1 -296
rect 16 -302 18 -296
rect 49 -297 52 -296
rect 5 -311 7 -305
rect 23 -311 25 -304
rect 57 -306 60 -301
rect 41 -310 51 -307
rect 57 -309 63 -306
rect 41 -311 43 -310
rect 5 -313 43 -311
rect 57 -311 60 -309
rect 23 -317 25 -313
rect 49 -318 52 -315
rect -1 -322 1 -320
rect 49 -320 60 -318
rect 49 -322 53 -320
rect -13 -324 53 -322
<< labels >>
rlabel polysilicon 21 59 21 59 1 a3
rlabel polysilicon 21 5 21 5 1 a2
rlabel polysilicon 21 -41 21 -41 1 a1
rlabel polysilicon 21 -100 21 -100 1 a0
rlabel metal1 60 -93 60 -93 1 and_a0
rlabel metal1 60 -34 60 -34 1 and_a1
rlabel metal1 60 12 60 12 1 and_a2
rlabel metal1 61 68 61 68 1 and_a3
rlabel polysilicon -16 56 -16 56 1 D3
rlabel metal1 28 80 28 80 1 vdd
rlabel metal1 36 52 36 52 1 gnd
rlabel polysilicon 21 -154 21 -154 1 b3
rlabel polysilicon 21 -210 21 -210 1 b2
rlabel polysilicon 21 -256 21 -256 1 b1
rlabel polysilicon 21 -315 21 -315 1 b0
rlabel metal1 60 -308 60 -308 1 and_b0
rlabel metal1 61 -249 61 -249 1 and_b1
rlabel metal1 62 -203 62 -203 1 and_b2
rlabel metal1 61 -148 61 -148 1 and_b3
<< end >>
