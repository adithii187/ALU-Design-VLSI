magic
tech scmos
timestamp 1701523314
<< nwell >>
rect -30258 9675 -30150 10350
rect -29448 9675 -29340 10350
rect -28566 9675 -28458 10350
rect -28908 9486 -28719 9540
rect -29934 9423 -29745 9477
rect -30402 9270 -30078 9360
rect -29934 9315 -29781 9423
rect -29376 9333 -29052 9423
rect -28908 9378 -28755 9486
rect -28908 9369 -28845 9378
rect -28827 9369 -28755 9378
rect -29934 9306 -29871 9315
rect -29853 9306 -29781 9315
rect -29718 8919 -29367 9036
rect -30258 7578 -30150 8253
rect -29448 7578 -29340 8253
rect -28566 7578 -28458 8253
rect -28908 7389 -28719 7443
rect -29934 7326 -29745 7380
rect -30402 7173 -30078 7263
rect -29934 7218 -29781 7326
rect -29376 7236 -29052 7326
rect -28908 7281 -28755 7389
rect -28908 7272 -28845 7281
rect -28827 7272 -28755 7281
rect -29934 7209 -29871 7218
rect -29853 7209 -29781 7218
rect -29718 6822 -29367 6939
rect -30258 5463 -30150 6138
rect -29448 5463 -29340 6138
rect -28566 5463 -28458 6138
rect -28908 5274 -28719 5328
rect -29934 5211 -29745 5265
rect -30402 5058 -30078 5148
rect -29934 5103 -29781 5211
rect -29376 5121 -29052 5211
rect -28908 5166 -28755 5274
rect -28908 5157 -28845 5166
rect -28827 5157 -28755 5166
rect -29934 5094 -29871 5103
rect -29853 5094 -29781 5103
rect -29718 4707 -29367 4824
rect -30258 3528 -30150 4203
rect -29448 3528 -29340 4203
rect -28566 3528 -28458 4203
rect -28908 3339 -28719 3393
rect -29934 3276 -29745 3330
rect -30402 3123 -30078 3213
rect -29934 3168 -29781 3276
rect -29376 3186 -29052 3276
rect -28908 3231 -28755 3339
rect -28908 3222 -28845 3231
rect -28827 3222 -28755 3231
rect -29934 3159 -29871 3168
rect -29853 3159 -29781 3168
rect -29718 2772 -29367 2889
rect -29898 -162 -29790 513
rect -29547 441 -29358 486
rect -29538 333 -29385 441
rect -29538 324 -29475 333
rect -29457 324 -29385 333
rect -29178 135 -28989 180
rect -28332 171 -28143 225
rect -29169 27 -29016 135
rect -29169 18 -29106 27
rect -29088 18 -29016 27
rect -28800 18 -28476 108
rect -28332 63 -28179 171
rect -28332 54 -28269 63
rect -28251 54 -28179 63
rect -33462 -243 -33273 -189
rect -33930 -396 -33606 -306
rect -33462 -351 -33309 -243
rect -33462 -360 -33399 -351
rect -33381 -360 -33309 -351
rect -33462 -738 -33273 -684
rect -33930 -891 -33606 -801
rect -33462 -846 -33309 -738
rect -33462 -855 -33399 -846
rect -33381 -855 -33309 -846
rect -34488 -1134 -34137 -1017
rect -33462 -1152 -33273 -1098
rect -29898 -1107 -29790 -432
rect -29547 -504 -29358 -459
rect -29538 -612 -29385 -504
rect -29538 -621 -29475 -612
rect -29457 -621 -29385 -612
rect -29196 -657 -29007 -630
rect -29205 -675 -29007 -657
rect -28404 -639 -28215 -585
rect -27576 -639 -27387 -585
rect -29187 -783 -29034 -675
rect -29187 -792 -29124 -783
rect -29106 -792 -29034 -783
rect -28872 -792 -28548 -702
rect -28404 -747 -28251 -639
rect -28404 -756 -28341 -747
rect -28323 -756 -28251 -747
rect -28044 -792 -27720 -702
rect -27576 -747 -27423 -639
rect -27126 -675 -27108 -666
rect -27576 -756 -27513 -747
rect -27495 -756 -27423 -747
rect -27144 -792 -26622 -675
rect -26838 -810 -26802 -792
rect -33930 -1305 -33606 -1215
rect -33462 -1260 -33309 -1152
rect -33462 -1269 -33399 -1260
rect -33381 -1269 -33309 -1260
rect -28728 -1431 -27738 -1404
rect -33462 -1683 -33273 -1629
rect -33930 -1836 -33606 -1746
rect -33462 -1791 -33309 -1683
rect -33462 -1800 -33399 -1791
rect -33381 -1800 -33309 -1791
rect -29898 -2124 -29790 -1449
rect -28737 -1458 -27738 -1431
rect -29547 -1521 -29367 -1476
rect -29214 -1521 -29025 -1476
rect -29538 -1629 -29385 -1521
rect -29538 -1638 -29475 -1629
rect -29457 -1638 -29385 -1629
rect -29205 -1629 -29052 -1521
rect -28728 -1566 -27738 -1458
rect -29205 -1638 -29142 -1629
rect -29124 -1638 -29052 -1629
rect -33462 -2250 -33273 -2196
rect -33930 -2403 -33606 -2313
rect -33462 -2358 -33309 -2250
rect -33462 -2367 -33399 -2358
rect -33381 -2367 -33309 -2358
rect -33462 -2745 -33273 -2691
rect -28881 -2727 -27891 -2700
rect -33930 -2898 -33606 -2808
rect -33462 -2853 -33309 -2745
rect -33462 -2862 -33399 -2853
rect -33381 -2862 -33309 -2853
rect -33462 -3159 -33273 -3105
rect -33930 -3312 -33606 -3222
rect -33462 -3267 -33309 -3159
rect -33462 -3276 -33399 -3267
rect -33381 -3276 -33309 -3267
rect -29898 -3420 -29790 -2745
rect -28890 -2754 -27891 -2727
rect -29547 -2817 -29367 -2772
rect -29268 -2817 -29079 -2772
rect -29538 -2925 -29385 -2817
rect -29538 -2934 -29475 -2925
rect -29457 -2934 -29385 -2925
rect -29259 -2925 -29106 -2817
rect -28881 -2862 -27891 -2754
rect -29259 -2934 -29196 -2925
rect -29178 -2934 -29106 -2925
rect -33462 -3690 -33273 -3636
rect -33930 -3843 -33606 -3753
rect -33462 -3798 -33309 -3690
rect -33462 -3807 -33399 -3798
rect -33381 -3807 -33309 -3798
rect -29898 -4491 -29790 -3816
rect -29547 -3888 -29358 -3843
rect -29538 -3996 -29385 -3888
rect -29538 -4005 -29475 -3996
rect -29457 -4005 -29385 -3996
rect -29178 -4194 -28989 -4149
rect -28332 -4158 -28143 -4104
rect -29169 -4302 -29016 -4194
rect -29169 -4311 -29106 -4302
rect -29088 -4311 -29016 -4302
rect -28800 -4311 -28476 -4221
rect -28332 -4266 -28179 -4158
rect -28332 -4275 -28269 -4266
rect -28251 -4275 -28179 -4266
rect -29898 -5436 -29790 -4761
rect -29547 -4833 -29358 -4788
rect -29538 -4941 -29385 -4833
rect -29538 -4950 -29475 -4941
rect -29457 -4950 -29385 -4941
rect -29196 -4986 -29007 -4959
rect -29205 -5004 -29007 -4986
rect -28404 -4968 -28215 -4914
rect -27576 -4941 -27387 -4914
rect -27576 -4959 -27108 -4941
rect -27576 -4968 -27387 -4959
rect -29187 -5112 -29034 -5004
rect -29187 -5121 -29124 -5112
rect -29106 -5121 -29034 -5112
rect -28872 -5121 -28548 -5031
rect -28404 -5076 -28251 -4968
rect -28404 -5085 -28341 -5076
rect -28323 -5085 -28251 -5076
rect -28044 -5121 -27720 -5031
rect -27576 -5076 -27423 -4968
rect -27126 -5004 -27108 -4959
rect -27576 -5085 -27513 -5076
rect -27495 -5085 -27423 -5076
rect -27144 -5121 -26622 -5004
rect -26838 -5139 -26802 -5121
rect -28728 -5760 -27738 -5733
rect -29898 -6453 -29790 -5778
rect -28737 -5787 -27738 -5760
rect -29547 -5850 -29367 -5805
rect -29214 -5850 -29025 -5805
rect -29538 -5958 -29385 -5850
rect -29538 -5967 -29475 -5958
rect -29457 -5967 -29385 -5958
rect -29205 -5958 -29052 -5850
rect -28728 -5895 -27738 -5787
rect -29205 -5967 -29142 -5958
rect -29124 -5967 -29052 -5958
rect -28881 -7056 -27891 -7029
rect -29898 -7749 -29790 -7074
rect -28890 -7083 -27891 -7056
rect -29547 -7146 -29367 -7101
rect -29268 -7146 -29079 -7101
rect -29538 -7254 -29385 -7146
rect -29538 -7263 -29475 -7254
rect -29457 -7263 -29385 -7254
rect -29259 -7254 -29106 -7146
rect -28881 -7191 -27891 -7083
rect -29259 -7263 -29196 -7254
rect -29178 -7263 -29106 -7254
rect -33444 -8100 -33255 -8046
rect -33912 -8253 -33588 -8163
rect -33444 -8208 -33291 -8100
rect -33444 -8217 -33381 -8208
rect -33363 -8217 -33291 -8208
rect -33444 -8595 -33255 -8541
rect -33912 -8748 -33588 -8658
rect -33444 -8703 -33291 -8595
rect -33444 -8712 -33381 -8703
rect -33363 -8712 -33291 -8703
rect -33444 -9009 -33255 -8955
rect -33912 -9162 -33588 -9072
rect -33444 -9117 -33291 -9009
rect -33444 -9126 -33381 -9117
rect -33363 -9126 -33291 -9117
rect -29898 -9288 -29790 -8613
rect -29547 -8685 -29358 -8640
rect -29538 -8793 -29385 -8685
rect -29538 -8802 -29475 -8793
rect -29457 -8802 -29385 -8793
rect -33444 -9540 -33255 -9486
rect -33912 -9693 -33588 -9603
rect -33444 -9648 -33291 -9540
rect -33444 -9657 -33381 -9648
rect -33363 -9657 -33291 -9648
rect -33444 -10017 -33255 -9963
rect -33912 -10170 -33588 -10080
rect -33444 -10125 -33291 -10017
rect -33444 -10134 -33381 -10125
rect -33363 -10134 -33291 -10125
rect -29898 -10233 -29790 -9558
rect -29547 -9630 -29358 -9585
rect -29538 -9738 -29385 -9630
rect -29538 -9747 -29475 -9738
rect -29457 -9747 -29385 -9738
rect -28260 -9846 -27270 -9684
rect -26433 -9693 -26244 -9639
rect -26901 -9846 -26577 -9756
rect -26433 -9801 -26280 -9693
rect -26433 -9810 -26370 -9801
rect -26352 -9810 -26280 -9801
rect -33444 -10512 -33255 -10458
rect -33912 -10665 -33588 -10575
rect -33444 -10620 -33291 -10512
rect -33444 -10629 -33381 -10620
rect -33363 -10629 -33291 -10620
rect -33444 -10926 -33255 -10872
rect -33912 -11079 -33588 -10989
rect -33444 -11034 -33291 -10926
rect -33444 -11043 -33381 -11034
rect -33363 -11043 -33291 -11034
rect -29898 -11250 -29790 -10575
rect -29547 -10647 -29358 -10602
rect -29538 -10755 -29385 -10647
rect -29538 -10764 -29475 -10755
rect -29457 -10764 -29385 -10755
rect -35442 -11439 -35253 -11385
rect -35910 -11592 -35586 -11502
rect -35442 -11547 -35289 -11439
rect -33444 -11457 -33255 -11403
rect -35442 -11556 -35379 -11547
rect -35361 -11556 -35289 -11547
rect -33912 -11610 -33588 -11520
rect -33444 -11565 -33291 -11457
rect -33444 -11574 -33381 -11565
rect -33363 -11574 -33291 -11565
rect -35442 -11907 -35253 -11853
rect -36243 -12078 -36054 -12051
rect -35910 -12060 -35586 -11970
rect -35442 -12015 -35289 -11907
rect -35442 -12024 -35379 -12015
rect -35361 -12024 -35289 -12015
rect -36243 -12096 -36216 -12078
rect -36108 -12096 -36054 -12078
rect -36234 -12204 -36081 -12096
rect -36234 -12213 -36171 -12204
rect -36153 -12213 -36081 -12204
rect -35442 -12348 -35253 -12294
rect -33444 -12321 -33255 -12267
rect -36234 -12393 -36045 -12375
rect -35973 -12393 -35955 -12366
rect -36234 -12411 -35955 -12393
rect -36234 -12420 -36045 -12411
rect -36225 -12528 -36072 -12420
rect -35910 -12501 -35586 -12411
rect -35442 -12456 -35289 -12348
rect -35442 -12465 -35379 -12456
rect -35361 -12465 -35289 -12456
rect -33912 -12474 -33588 -12384
rect -33444 -12429 -33291 -12321
rect -33444 -12438 -33381 -12429
rect -33363 -12438 -33291 -12429
rect -36225 -12537 -36162 -12528
rect -36144 -12537 -36072 -12528
rect -29898 -12546 -29790 -11871
rect -29547 -11916 -29358 -11898
rect -29547 -11934 -29349 -11916
rect -29547 -11943 -29358 -11934
rect -29538 -12051 -29385 -11943
rect -29538 -12060 -29475 -12051
rect -29457 -12060 -29385 -12051
rect -35442 -12762 -35253 -12708
rect -35910 -12915 -35586 -12825
rect -35442 -12870 -35289 -12762
rect -35442 -12879 -35379 -12870
rect -35361 -12879 -35289 -12870
rect -33444 -12816 -33255 -12762
rect -33912 -12969 -33588 -12879
rect -33444 -12924 -33291 -12816
rect -33444 -12933 -33381 -12924
rect -33363 -12933 -33291 -12924
rect -33444 -13230 -33255 -13176
rect -33912 -13383 -33588 -13293
rect -33444 -13338 -33291 -13230
rect -33444 -13347 -33381 -13338
rect -33363 -13347 -33291 -13338
rect -33444 -13761 -33255 -13707
rect -33912 -13914 -33588 -13824
rect -33444 -13869 -33291 -13761
rect -31473 -13770 -31284 -13716
rect -33444 -13878 -33381 -13869
rect -33363 -13878 -33291 -13869
rect -31941 -13923 -31617 -13833
rect -31473 -13878 -31320 -13770
rect -31473 -13887 -31410 -13878
rect -31392 -13887 -31320 -13878
rect -33444 -14256 -33255 -14202
rect -31473 -14247 -31284 -14193
rect -33912 -14409 -33588 -14319
rect -33444 -14364 -33291 -14256
rect -33444 -14373 -33381 -14364
rect -33363 -14373 -33291 -14364
rect -31941 -14400 -31617 -14310
rect -31473 -14355 -31320 -14247
rect -31473 -14364 -31410 -14355
rect -31392 -14364 -31320 -14355
rect -31473 -14643 -31284 -14589
rect -33444 -14751 -33255 -14697
rect -33912 -14904 -33588 -14814
rect -33444 -14859 -33291 -14751
rect -31941 -14796 -31617 -14706
rect -31473 -14751 -31320 -14643
rect -31473 -14760 -31410 -14751
rect -31392 -14760 -31320 -14751
rect -33444 -14868 -33381 -14859
rect -33363 -14868 -33291 -14859
rect -31473 -15111 -31284 -15057
rect -33444 -15165 -33255 -15111
rect -33912 -15318 -33588 -15228
rect -33444 -15273 -33291 -15165
rect -31941 -15264 -31617 -15174
rect -31473 -15219 -31320 -15111
rect -31473 -15228 -31410 -15219
rect -31392 -15228 -31320 -15219
rect -33444 -15282 -33381 -15273
rect -33363 -15282 -33291 -15273
rect -33444 -15696 -33255 -15642
rect -33912 -15849 -33588 -15759
rect -33444 -15804 -33291 -15696
rect -33444 -15813 -33381 -15804
rect -33363 -15813 -33291 -15804
<< ntransistor >>
rect -30483 10269 -30429 10287
rect -29673 10269 -29619 10287
rect -30483 10098 -30429 10116
rect -30483 9900 -30429 9918
rect -30483 9738 -30429 9756
rect -28791 10269 -28737 10287
rect -29673 10098 -29619 10116
rect -29673 9900 -29619 9918
rect -29673 9738 -29619 9756
rect -28791 10098 -28737 10116
rect -28791 9900 -28737 9918
rect -28791 9738 -28737 9756
rect -29871 9225 -29853 9252
rect -30330 9171 -30312 9198
rect -30168 9171 -30150 9198
rect -29304 9234 -29286 9261
rect -29142 9234 -29124 9261
rect -28845 9288 -28827 9315
rect -29655 8820 -29637 8847
rect -29565 8820 -29547 8847
rect -29439 8820 -29421 8847
rect -30483 8172 -30429 8190
rect -29673 8172 -29619 8190
rect -30483 8001 -30429 8019
rect -30483 7803 -30429 7821
rect -30483 7641 -30429 7659
rect -28791 8172 -28737 8190
rect -29673 8001 -29619 8019
rect -29673 7803 -29619 7821
rect -29673 7641 -29619 7659
rect -28791 8001 -28737 8019
rect -28791 7803 -28737 7821
rect -28791 7641 -28737 7659
rect -29871 7128 -29853 7155
rect -30330 7074 -30312 7101
rect -30168 7074 -30150 7101
rect -29304 7137 -29286 7164
rect -29142 7137 -29124 7164
rect -28845 7191 -28827 7218
rect -29655 6723 -29637 6750
rect -29565 6723 -29547 6750
rect -29439 6723 -29421 6750
rect -30483 6057 -30429 6075
rect -29673 6057 -29619 6075
rect -30483 5886 -30429 5904
rect -30483 5688 -30429 5706
rect -30483 5526 -30429 5544
rect -28791 6057 -28737 6075
rect -29673 5886 -29619 5904
rect -29673 5688 -29619 5706
rect -29673 5526 -29619 5544
rect -28791 5886 -28737 5904
rect -28791 5688 -28737 5706
rect -28791 5526 -28737 5544
rect -29871 5013 -29853 5040
rect -30330 4959 -30312 4986
rect -30168 4959 -30150 4986
rect -29304 5022 -29286 5049
rect -29142 5022 -29124 5049
rect -28845 5076 -28827 5103
rect -29655 4608 -29637 4635
rect -29565 4608 -29547 4635
rect -29439 4608 -29421 4635
rect -30483 4122 -30429 4140
rect -29673 4122 -29619 4140
rect -30483 3951 -30429 3969
rect -30483 3753 -30429 3771
rect -30483 3591 -30429 3609
rect -28791 4122 -28737 4140
rect -29673 3951 -29619 3969
rect -29673 3753 -29619 3771
rect -29673 3591 -29619 3609
rect -28791 3951 -28737 3969
rect -28791 3753 -28737 3771
rect -28791 3591 -28737 3609
rect -29871 3078 -29853 3105
rect -30330 3024 -30312 3051
rect -30168 3024 -30150 3051
rect -29304 3087 -29286 3114
rect -29142 3087 -29124 3114
rect -28845 3141 -28827 3168
rect -29655 2673 -29637 2700
rect -29565 2673 -29547 2700
rect -29439 2673 -29421 2700
rect -30123 432 -30069 450
rect -30123 261 -30069 279
rect -29475 243 -29457 270
rect -30123 63 -30069 81
rect -30123 -99 -30069 -81
rect -29106 -63 -29088 -36
rect -28269 -27 -28251 0
rect -28728 -81 -28710 -54
rect -28620 -81 -28611 -54
rect -28566 -81 -28548 -54
rect -33399 -441 -33381 -414
rect -33858 -495 -33840 -468
rect -33696 -495 -33678 -468
rect -30123 -513 -30069 -495
rect -33399 -936 -33381 -909
rect -33858 -990 -33840 -963
rect -33696 -990 -33678 -963
rect -34425 -1233 -34407 -1206
rect -34335 -1233 -34317 -1206
rect -34209 -1233 -34191 -1206
rect -33399 -1350 -33381 -1323
rect -33858 -1404 -33840 -1377
rect -33696 -1404 -33678 -1377
rect -33399 -1881 -33381 -1854
rect -33858 -1935 -33840 -1908
rect -33696 -1935 -33678 -1908
rect -33399 -2448 -33381 -2421
rect -33858 -2502 -33840 -2475
rect -33696 -2502 -33678 -2475
rect -33399 -2943 -33381 -2916
rect -33858 -2997 -33840 -2970
rect -33696 -2997 -33678 -2970
rect -33399 -3357 -33381 -3330
rect -33858 -3411 -33840 -3384
rect -33696 -3411 -33678 -3384
rect -33399 -3888 -33381 -3861
rect -33858 -3942 -33840 -3915
rect -33696 -3942 -33678 -3915
rect -30123 -684 -30069 -666
rect -29475 -702 -29457 -675
rect -30123 -882 -30069 -864
rect -29124 -873 -29106 -846
rect -28341 -837 -28323 -810
rect -27513 -837 -27495 -810
rect -28800 -891 -28782 -864
rect -28692 -891 -28683 -864
rect -28638 -891 -28620 -864
rect -27972 -891 -27954 -864
rect -27810 -891 -27792 -864
rect -27090 -891 -27072 -864
rect -27000 -891 -26982 -864
rect -26910 -891 -26892 -864
rect -26820 -891 -26802 -864
rect -26694 -891 -26676 -864
rect -30123 -1044 -30069 -1026
rect -30123 -1530 -30069 -1512
rect -30123 -1701 -30069 -1683
rect -29475 -1719 -29457 -1692
rect -29142 -1719 -29124 -1692
rect -28638 -1701 -28620 -1674
rect -28512 -1701 -28494 -1674
rect -28368 -1701 -28350 -1674
rect -28242 -1701 -28224 -1674
rect -28107 -1701 -28089 -1674
rect -27846 -1701 -27828 -1674
rect -30123 -1899 -30069 -1881
rect -30123 -2061 -30069 -2043
rect -30123 -2826 -30069 -2808
rect -30123 -2997 -30069 -2979
rect -29475 -3015 -29457 -2988
rect -29196 -3015 -29178 -2988
rect -28791 -2997 -28773 -2970
rect -28665 -2997 -28647 -2970
rect -28521 -2997 -28503 -2970
rect -28395 -2997 -28377 -2970
rect -28260 -2997 -28242 -2970
rect -27999 -2997 -27981 -2970
rect -30123 -3195 -30069 -3177
rect -30123 -3357 -30069 -3339
rect -30123 -3897 -30069 -3879
rect -30123 -4068 -30069 -4050
rect -29475 -4086 -29457 -4059
rect -30123 -4266 -30069 -4248
rect -30123 -4428 -30069 -4410
rect -29106 -4392 -29088 -4365
rect -28269 -4356 -28251 -4329
rect -28728 -4410 -28710 -4383
rect -28620 -4410 -28611 -4383
rect -28566 -4410 -28548 -4383
rect -30123 -4842 -30069 -4824
rect -30123 -5013 -30069 -4995
rect -29475 -5031 -29457 -5004
rect -30123 -5211 -30069 -5193
rect -29124 -5202 -29106 -5175
rect -28341 -5166 -28323 -5139
rect -27513 -5166 -27495 -5139
rect -28800 -5220 -28782 -5193
rect -28692 -5220 -28683 -5193
rect -28638 -5220 -28620 -5193
rect -27972 -5220 -27954 -5193
rect -27810 -5220 -27792 -5193
rect -27090 -5220 -27072 -5193
rect -27000 -5220 -26982 -5193
rect -26910 -5220 -26892 -5193
rect -26820 -5220 -26802 -5193
rect -26694 -5220 -26676 -5193
rect -30123 -5373 -30069 -5355
rect -30123 -5859 -30069 -5841
rect -30123 -6030 -30069 -6012
rect -29475 -6048 -29457 -6021
rect -29142 -6048 -29124 -6021
rect -28638 -6030 -28620 -6003
rect -28512 -6030 -28494 -6003
rect -28368 -6030 -28350 -6003
rect -28242 -6030 -28224 -6003
rect -28107 -6030 -28089 -6003
rect -27846 -6030 -27828 -6003
rect -30123 -6228 -30069 -6210
rect -30123 -6390 -30069 -6372
rect -33381 -8298 -33363 -8271
rect -33840 -8352 -33822 -8325
rect -33678 -8352 -33660 -8325
rect -33381 -8793 -33363 -8766
rect -33840 -8847 -33822 -8820
rect -33678 -8847 -33660 -8820
rect -33381 -9207 -33363 -9180
rect -33840 -9261 -33822 -9234
rect -33678 -9261 -33660 -9234
rect -33381 -9738 -33363 -9711
rect -33840 -9792 -33822 -9765
rect -33678 -9792 -33660 -9765
rect -33381 -10215 -33363 -10188
rect -33840 -10269 -33822 -10242
rect -33678 -10269 -33660 -10242
rect -35379 -11637 -35361 -11610
rect -35838 -11691 -35820 -11664
rect -35676 -11691 -35658 -11664
rect -33381 -10710 -33363 -10683
rect -33840 -10764 -33822 -10737
rect -33678 -10764 -33660 -10737
rect -33381 -11124 -33363 -11097
rect -33840 -11178 -33822 -11151
rect -33678 -11178 -33660 -11151
rect -30123 -7155 -30069 -7137
rect -30123 -7326 -30069 -7308
rect -29475 -7344 -29457 -7317
rect -30123 -7524 -30069 -7506
rect -30123 -7686 -30069 -7668
rect -30123 -8694 -30069 -8676
rect -29196 -7344 -29178 -7317
rect -28791 -7326 -28773 -7299
rect -28665 -7326 -28647 -7299
rect -28521 -7326 -28503 -7299
rect -28395 -7326 -28377 -7299
rect -28260 -7326 -28242 -7299
rect -27999 -7326 -27981 -7299
rect -30123 -8865 -30069 -8847
rect -29475 -8883 -29457 -8856
rect -30123 -9063 -30069 -9045
rect -30123 -9225 -30069 -9207
rect -30123 -9639 -30069 -9621
rect -30123 -9810 -30069 -9792
rect -29475 -9828 -29457 -9801
rect -30123 -10008 -30069 -9990
rect -26370 -9891 -26352 -9864
rect -26829 -9945 -26811 -9918
rect -26667 -9945 -26649 -9918
rect -28170 -9981 -28152 -9954
rect -28044 -9981 -28026 -9954
rect -27900 -9981 -27882 -9954
rect -27774 -9981 -27756 -9954
rect -27639 -9981 -27621 -9954
rect -27378 -9981 -27360 -9954
rect -30123 -10170 -30069 -10152
rect -30123 -10656 -30069 -10638
rect -30123 -10827 -30069 -10809
rect -29475 -10845 -29457 -10818
rect -30123 -11025 -30069 -11007
rect -30123 -11187 -30069 -11169
rect -35379 -12105 -35361 -12078
rect -35838 -12159 -35820 -12132
rect -35676 -12159 -35658 -12132
rect -36171 -12294 -36153 -12267
rect -33381 -11655 -33363 -11628
rect -33840 -11709 -33822 -11682
rect -33678 -11709 -33660 -11682
rect -30123 -11952 -30069 -11934
rect -35379 -12546 -35361 -12519
rect -36162 -12618 -36144 -12591
rect -35838 -12600 -35820 -12573
rect -35703 -12600 -35685 -12573
rect -35676 -12600 -35658 -12573
rect -33381 -12519 -33363 -12492
rect -33840 -12573 -33822 -12546
rect -33678 -12573 -33660 -12546
rect -30123 -12123 -30069 -12105
rect -29475 -12141 -29457 -12114
rect -30123 -12321 -30069 -12303
rect -30123 -12483 -30069 -12465
rect -35379 -12960 -35361 -12933
rect -35838 -13014 -35820 -12987
rect -35721 -13014 -35703 -12987
rect -35676 -13014 -35658 -12987
rect -33381 -13014 -33363 -12987
rect -33840 -13068 -33822 -13041
rect -33678 -13068 -33660 -13041
rect -33381 -13428 -33363 -13401
rect -33840 -13482 -33822 -13455
rect -33678 -13482 -33660 -13455
rect -33381 -13959 -33363 -13932
rect -33840 -14013 -33822 -13986
rect -33678 -14013 -33660 -13986
rect -31410 -13968 -31392 -13941
rect -31869 -14022 -31851 -13995
rect -31707 -14022 -31689 -13995
rect -33381 -14454 -33363 -14427
rect -31410 -14445 -31392 -14418
rect -33840 -14508 -33822 -14481
rect -33678 -14508 -33660 -14481
rect -31869 -14499 -31851 -14472
rect -31707 -14499 -31689 -14472
rect -31410 -14841 -31392 -14814
rect -31869 -14895 -31851 -14868
rect -31707 -14895 -31689 -14868
rect -33381 -14949 -33363 -14922
rect -33840 -15003 -33822 -14976
rect -33678 -15003 -33660 -14976
rect -31410 -15309 -31392 -15282
rect -33381 -15363 -33363 -15336
rect -31869 -15363 -31851 -15336
rect -31707 -15363 -31689 -15336
rect -33840 -15417 -33822 -15390
rect -33678 -15417 -33660 -15390
rect -33381 -15894 -33363 -15867
rect -33840 -15948 -33822 -15921
rect -33678 -15948 -33660 -15921
<< ptransistor >>
rect -30231 10269 -30168 10287
rect -29421 10269 -29358 10287
rect -30231 10098 -30168 10116
rect -30231 9900 -30168 9918
rect -30231 9738 -30168 9756
rect -28539 10269 -28476 10287
rect -29421 10098 -29358 10116
rect -29421 9900 -29358 9918
rect -29421 9738 -29358 9756
rect -28539 10098 -28476 10116
rect -28539 9900 -28476 9918
rect -28539 9738 -28476 9756
rect -30330 9297 -30312 9342
rect -30168 9297 -30150 9342
rect -29871 9324 -29853 9378
rect -29304 9360 -29286 9405
rect -29142 9360 -29124 9405
rect -28845 9387 -28827 9441
rect -29655 8937 -29637 8982
rect -29565 8937 -29547 8982
rect -29439 8937 -29421 8982
rect -30231 8172 -30168 8190
rect -29421 8172 -29358 8190
rect -30231 8001 -30168 8019
rect -30231 7803 -30168 7821
rect -30231 7641 -30168 7659
rect -28539 8172 -28476 8190
rect -29421 8001 -29358 8019
rect -29421 7803 -29358 7821
rect -29421 7641 -29358 7659
rect -28539 8001 -28476 8019
rect -28539 7803 -28476 7821
rect -28539 7641 -28476 7659
rect -30330 7200 -30312 7245
rect -30168 7200 -30150 7245
rect -29871 7227 -29853 7281
rect -29304 7263 -29286 7308
rect -29142 7263 -29124 7308
rect -28845 7290 -28827 7344
rect -29655 6840 -29637 6885
rect -29565 6840 -29547 6885
rect -29439 6840 -29421 6885
rect -30231 6057 -30168 6075
rect -29421 6057 -29358 6075
rect -30231 5886 -30168 5904
rect -30231 5688 -30168 5706
rect -30231 5526 -30168 5544
rect -28539 6057 -28476 6075
rect -29421 5886 -29358 5904
rect -29421 5688 -29358 5706
rect -29421 5526 -29358 5544
rect -28539 5886 -28476 5904
rect -28539 5688 -28476 5706
rect -28539 5526 -28476 5544
rect -30330 5085 -30312 5130
rect -30168 5085 -30150 5130
rect -29871 5112 -29853 5166
rect -29304 5148 -29286 5193
rect -29142 5148 -29124 5193
rect -28845 5175 -28827 5229
rect -29655 4725 -29637 4770
rect -29565 4725 -29547 4770
rect -29439 4725 -29421 4770
rect -30231 4122 -30168 4140
rect -29421 4122 -29358 4140
rect -30231 3951 -30168 3969
rect -30231 3753 -30168 3771
rect -30231 3591 -30168 3609
rect -28539 4122 -28476 4140
rect -29421 3951 -29358 3969
rect -29421 3753 -29358 3771
rect -29421 3591 -29358 3609
rect -28539 3951 -28476 3969
rect -28539 3753 -28476 3771
rect -28539 3591 -28476 3609
rect -30330 3150 -30312 3195
rect -30168 3150 -30150 3195
rect -29871 3177 -29853 3231
rect -29304 3213 -29286 3258
rect -29142 3213 -29124 3258
rect -28845 3240 -28827 3294
rect -29655 2790 -29637 2835
rect -29565 2790 -29547 2835
rect -29439 2790 -29421 2835
rect -29871 432 -29808 450
rect -29475 342 -29457 396
rect -29871 261 -29808 279
rect -29871 63 -29808 81
rect -29871 -99 -29808 -81
rect -29106 36 -29088 90
rect -28728 45 -28710 90
rect -28566 45 -28548 90
rect -28269 72 -28251 126
rect -33858 -369 -33840 -324
rect -33696 -369 -33678 -324
rect -33399 -342 -33381 -288
rect -29871 -513 -29808 -495
rect -33858 -864 -33840 -819
rect -33696 -864 -33678 -819
rect -33399 -837 -33381 -783
rect -34425 -1116 -34407 -1071
rect -34335 -1116 -34317 -1071
rect -34209 -1116 -34191 -1071
rect -33858 -1278 -33840 -1233
rect -33696 -1278 -33678 -1233
rect -33399 -1251 -33381 -1197
rect -33858 -1809 -33840 -1764
rect -33696 -1809 -33678 -1764
rect -33399 -1782 -33381 -1728
rect -33858 -2376 -33840 -2331
rect -33696 -2376 -33678 -2331
rect -33399 -2349 -33381 -2295
rect -33858 -2871 -33840 -2826
rect -33696 -2871 -33678 -2826
rect -33399 -2844 -33381 -2790
rect -33858 -3285 -33840 -3240
rect -33696 -3285 -33678 -3240
rect -33399 -3258 -33381 -3204
rect -33858 -3816 -33840 -3771
rect -33696 -3816 -33678 -3771
rect -33399 -3789 -33381 -3735
rect -33840 -8226 -33822 -8181
rect -33678 -8226 -33660 -8181
rect -33381 -8199 -33363 -8145
rect -29475 -603 -29457 -549
rect -29871 -684 -29808 -666
rect -29871 -882 -29808 -864
rect -29124 -774 -29106 -720
rect -28800 -765 -28782 -720
rect -28638 -765 -28620 -720
rect -28341 -738 -28323 -684
rect -27972 -765 -27954 -720
rect -27810 -765 -27792 -720
rect -27513 -738 -27495 -684
rect -27090 -774 -27072 -729
rect -27036 -774 -27018 -729
rect -27000 -774 -26982 -729
rect -26910 -774 -26892 -729
rect -26820 -774 -26802 -729
rect -26694 -774 -26676 -729
rect -29871 -1044 -29808 -1026
rect -29871 -1530 -29808 -1512
rect -28638 -1548 -28620 -1494
rect -28512 -1548 -28494 -1494
rect -28368 -1548 -28350 -1494
rect -28242 -1548 -28224 -1494
rect -28107 -1548 -28089 -1494
rect -27846 -1548 -27828 -1494
rect -29475 -1620 -29457 -1566
rect -29142 -1620 -29124 -1566
rect -29871 -1701 -29808 -1683
rect -29871 -1899 -29808 -1881
rect -29871 -2061 -29808 -2043
rect -29871 -2826 -29808 -2808
rect -28791 -2844 -28773 -2790
rect -28665 -2844 -28647 -2790
rect -28521 -2844 -28503 -2790
rect -28395 -2844 -28377 -2790
rect -28260 -2844 -28242 -2790
rect -27999 -2844 -27981 -2790
rect -29475 -2916 -29457 -2862
rect -29196 -2916 -29178 -2862
rect -29871 -2997 -29808 -2979
rect -29871 -3195 -29808 -3177
rect -29871 -3357 -29808 -3339
rect -29871 -3897 -29808 -3879
rect -29475 -3987 -29457 -3933
rect -29871 -4068 -29808 -4050
rect -29871 -4266 -29808 -4248
rect -29871 -4428 -29808 -4410
rect -29106 -4293 -29088 -4239
rect -28728 -4284 -28710 -4239
rect -28566 -4284 -28548 -4239
rect -28269 -4257 -28251 -4203
rect -29871 -4842 -29808 -4824
rect -29475 -4932 -29457 -4878
rect -29871 -5013 -29808 -4995
rect -29871 -5211 -29808 -5193
rect -29124 -5103 -29106 -5049
rect -28800 -5094 -28782 -5049
rect -28638 -5094 -28620 -5049
rect -28341 -5067 -28323 -5013
rect -27972 -5094 -27954 -5049
rect -27810 -5094 -27792 -5049
rect -27513 -5067 -27495 -5013
rect -27090 -5103 -27072 -5058
rect -27036 -5103 -27018 -5058
rect -27000 -5103 -26982 -5058
rect -26910 -5103 -26892 -5058
rect -26820 -5103 -26802 -5058
rect -26694 -5103 -26676 -5058
rect -29871 -5373 -29808 -5355
rect -29871 -5859 -29808 -5841
rect -28638 -5877 -28620 -5823
rect -28512 -5877 -28494 -5823
rect -28368 -5877 -28350 -5823
rect -28242 -5877 -28224 -5823
rect -28107 -5877 -28089 -5823
rect -27846 -5877 -27828 -5823
rect -29475 -5949 -29457 -5895
rect -29142 -5949 -29124 -5895
rect -29871 -6030 -29808 -6012
rect -29871 -6228 -29808 -6210
rect -29871 -6390 -29808 -6372
rect -33840 -8721 -33822 -8676
rect -33678 -8721 -33660 -8676
rect -33381 -8694 -33363 -8640
rect -33840 -9135 -33822 -9090
rect -33678 -9135 -33660 -9090
rect -33381 -9108 -33363 -9054
rect -33840 -9666 -33822 -9621
rect -33678 -9666 -33660 -9621
rect -33381 -9639 -33363 -9585
rect -33840 -10143 -33822 -10098
rect -33678 -10143 -33660 -10098
rect -33381 -10116 -33363 -10062
rect -33840 -10638 -33822 -10593
rect -33678 -10638 -33660 -10593
rect -33381 -10611 -33363 -10557
rect -35838 -11565 -35820 -11520
rect -35676 -11565 -35658 -11520
rect -35379 -11538 -35361 -11484
rect -35838 -12033 -35820 -11988
rect -35676 -12033 -35658 -11988
rect -35379 -12006 -35361 -11952
rect -33840 -11052 -33822 -11007
rect -33678 -11052 -33660 -11007
rect -33381 -11025 -33363 -10971
rect -29871 -7155 -29808 -7137
rect -29475 -7245 -29457 -7191
rect -29871 -7326 -29808 -7308
rect -29871 -7524 -29808 -7506
rect -29871 -7686 -29808 -7668
rect -29871 -8694 -29808 -8676
rect -28791 -7173 -28773 -7119
rect -28665 -7173 -28647 -7119
rect -28521 -7173 -28503 -7119
rect -28395 -7173 -28377 -7119
rect -28260 -7173 -28242 -7119
rect -27999 -7173 -27981 -7119
rect -29196 -7245 -29178 -7191
rect -29475 -8784 -29457 -8730
rect -29871 -8865 -29808 -8847
rect -29871 -9063 -29808 -9045
rect -29871 -9225 -29808 -9207
rect -29871 -9639 -29808 -9621
rect -29475 -9729 -29457 -9675
rect -29871 -9810 -29808 -9792
rect -29871 -10008 -29808 -9990
rect -28170 -9828 -28152 -9774
rect -28044 -9828 -28026 -9774
rect -27900 -9828 -27882 -9774
rect -27774 -9828 -27756 -9774
rect -27639 -9828 -27621 -9774
rect -27378 -9828 -27360 -9774
rect -26829 -9819 -26811 -9774
rect -26667 -9819 -26649 -9774
rect -26370 -9792 -26352 -9738
rect -29871 -10170 -29808 -10152
rect -29871 -10656 -29808 -10638
rect -29475 -10746 -29457 -10692
rect -29871 -10827 -29808 -10809
rect -29871 -11025 -29808 -11007
rect -29871 -11187 -29808 -11169
rect -33840 -11583 -33822 -11538
rect -33678 -11583 -33660 -11538
rect -33381 -11556 -33363 -11502
rect -36171 -12195 -36153 -12141
rect -36162 -12519 -36144 -12465
rect -35838 -12474 -35820 -12429
rect -35676 -12474 -35658 -12429
rect -35379 -12447 -35361 -12393
rect -29871 -11952 -29808 -11934
rect -33840 -12447 -33822 -12402
rect -33678 -12447 -33660 -12402
rect -33381 -12420 -33363 -12366
rect -35838 -12888 -35820 -12843
rect -35676 -12888 -35658 -12843
rect -35379 -12861 -35361 -12807
rect -29475 -12042 -29457 -11988
rect -29871 -12123 -29808 -12105
rect -29871 -12321 -29808 -12303
rect -29871 -12483 -29808 -12465
rect -33840 -12942 -33822 -12897
rect -33678 -12942 -33660 -12897
rect -33381 -12915 -33363 -12861
rect -33840 -13356 -33822 -13311
rect -33678 -13356 -33660 -13311
rect -33381 -13329 -33363 -13275
rect -33840 -13887 -33822 -13842
rect -33678 -13887 -33660 -13842
rect -33381 -13860 -33363 -13806
rect -31869 -13896 -31851 -13851
rect -31707 -13896 -31689 -13851
rect -31410 -13869 -31392 -13815
rect -33840 -14382 -33822 -14337
rect -33678 -14382 -33660 -14337
rect -33381 -14355 -33363 -14301
rect -31869 -14373 -31851 -14328
rect -31707 -14373 -31689 -14328
rect -31410 -14346 -31392 -14292
rect -31869 -14769 -31851 -14724
rect -31707 -14769 -31689 -14724
rect -31410 -14742 -31392 -14688
rect -33840 -14877 -33822 -14832
rect -33678 -14877 -33660 -14832
rect -33381 -14850 -33363 -14796
rect -33840 -15291 -33822 -15246
rect -33678 -15291 -33660 -15246
rect -33381 -15264 -33363 -15210
rect -31869 -15237 -31851 -15192
rect -31707 -15237 -31689 -15192
rect -31410 -15210 -31392 -15156
rect -33840 -15822 -33822 -15777
rect -33678 -15822 -33660 -15777
rect -33381 -15795 -33363 -15741
<< ndiffusion >>
rect -30483 10332 -30429 10341
rect -30483 10296 -30474 10332
rect -30438 10296 -30429 10332
rect -30483 10287 -30429 10296
rect -30483 10260 -30429 10269
rect -30483 10224 -30474 10260
rect -30438 10224 -30429 10260
rect -30483 10215 -30429 10224
rect -30483 10161 -30429 10170
rect -30483 10125 -30474 10161
rect -30438 10125 -30429 10161
rect -30483 10116 -30429 10125
rect -29673 10332 -29619 10341
rect -29673 10296 -29664 10332
rect -29628 10296 -29619 10332
rect -29673 10287 -29619 10296
rect -30483 10089 -30429 10098
rect -30483 10053 -30474 10089
rect -30438 10053 -30429 10089
rect -30483 10044 -30429 10053
rect -30483 9972 -30429 9981
rect -30483 9936 -30474 9972
rect -30438 9936 -30429 9972
rect -30483 9918 -30429 9936
rect -30483 9891 -30429 9900
rect -30483 9855 -30474 9891
rect -30438 9855 -30429 9891
rect -30483 9846 -30429 9855
rect -30483 9810 -30429 9819
rect -30483 9774 -30474 9810
rect -30438 9774 -30429 9810
rect -30483 9756 -30429 9774
rect -30483 9729 -30429 9738
rect -30483 9693 -30474 9729
rect -30438 9693 -30429 9729
rect -30483 9684 -30429 9693
rect -29673 10260 -29619 10269
rect -29673 10224 -29664 10260
rect -29628 10224 -29619 10260
rect -29673 10215 -29619 10224
rect -29673 10161 -29619 10170
rect -29673 10125 -29664 10161
rect -29628 10125 -29619 10161
rect -29673 10116 -29619 10125
rect -28791 10332 -28737 10341
rect -28791 10296 -28782 10332
rect -28746 10296 -28737 10332
rect -28791 10287 -28737 10296
rect -29673 10089 -29619 10098
rect -29673 10053 -29664 10089
rect -29628 10053 -29619 10089
rect -29673 10044 -29619 10053
rect -29673 9972 -29619 9981
rect -29673 9936 -29664 9972
rect -29628 9936 -29619 9972
rect -29673 9918 -29619 9936
rect -29673 9891 -29619 9900
rect -29673 9855 -29664 9891
rect -29628 9855 -29619 9891
rect -29673 9846 -29619 9855
rect -29673 9810 -29619 9819
rect -29673 9774 -29664 9810
rect -29628 9774 -29619 9810
rect -29673 9756 -29619 9774
rect -29673 9729 -29619 9738
rect -29673 9693 -29664 9729
rect -29628 9693 -29619 9729
rect -29673 9684 -29619 9693
rect -28791 10260 -28737 10269
rect -28791 10224 -28782 10260
rect -28746 10224 -28737 10260
rect -28791 10215 -28737 10224
rect -28791 10161 -28737 10170
rect -28791 10125 -28782 10161
rect -28746 10125 -28737 10161
rect -28791 10116 -28737 10125
rect -28791 10089 -28737 10098
rect -28791 10053 -28782 10089
rect -28746 10053 -28737 10089
rect -28791 10044 -28737 10053
rect -28791 9972 -28737 9981
rect -28791 9936 -28782 9972
rect -28746 9936 -28737 9972
rect -28791 9918 -28737 9936
rect -28791 9891 -28737 9900
rect -28791 9855 -28782 9891
rect -28746 9855 -28737 9891
rect -28791 9846 -28737 9855
rect -28791 9810 -28737 9819
rect -28791 9774 -28782 9810
rect -28746 9774 -28737 9810
rect -28791 9756 -28737 9774
rect -28791 9729 -28737 9738
rect -28791 9693 -28782 9729
rect -28746 9693 -28737 9729
rect -28791 9684 -28737 9693
rect -29916 9243 -29871 9252
rect -29916 9225 -29907 9243
rect -29880 9225 -29871 9243
rect -29853 9225 -29835 9252
rect -29808 9225 -29799 9252
rect -30366 9189 -30330 9198
rect -30366 9171 -30357 9189
rect -30339 9171 -30330 9189
rect -30312 9171 -30168 9198
rect -30150 9180 -30141 9198
rect -30123 9180 -30114 9198
rect -30150 9171 -30114 9180
rect -29340 9252 -29304 9261
rect -29340 9234 -29331 9252
rect -29313 9234 -29304 9252
rect -29286 9234 -29142 9261
rect -29124 9243 -29115 9261
rect -29097 9243 -29088 9261
rect -29124 9234 -29088 9243
rect -28890 9306 -28845 9315
rect -28890 9288 -28881 9306
rect -28854 9288 -28845 9306
rect -28827 9288 -28809 9315
rect -28782 9288 -28773 9315
rect -29691 8829 -29682 8847
rect -29664 8829 -29655 8847
rect -29691 8820 -29655 8829
rect -29637 8829 -29628 8847
rect -29637 8820 -29610 8829
rect -29601 8829 -29592 8847
rect -29574 8829 -29565 8847
rect -29601 8820 -29565 8829
rect -29547 8829 -29538 8847
rect -29547 8820 -29520 8829
rect -29475 8829 -29466 8847
rect -29448 8829 -29439 8847
rect -29475 8820 -29439 8829
rect -29421 8829 -29412 8847
rect -29394 8829 -29385 8847
rect -29421 8820 -29385 8829
rect -30483 8235 -30429 8244
rect -30483 8199 -30474 8235
rect -30438 8199 -30429 8235
rect -30483 8190 -30429 8199
rect -30483 8163 -30429 8172
rect -30483 8127 -30474 8163
rect -30438 8127 -30429 8163
rect -30483 8118 -30429 8127
rect -30483 8064 -30429 8073
rect -30483 8028 -30474 8064
rect -30438 8028 -30429 8064
rect -30483 8019 -30429 8028
rect -29673 8235 -29619 8244
rect -29673 8199 -29664 8235
rect -29628 8199 -29619 8235
rect -29673 8190 -29619 8199
rect -30483 7992 -30429 8001
rect -30483 7956 -30474 7992
rect -30438 7956 -30429 7992
rect -30483 7947 -30429 7956
rect -30483 7875 -30429 7884
rect -30483 7839 -30474 7875
rect -30438 7839 -30429 7875
rect -30483 7821 -30429 7839
rect -30483 7794 -30429 7803
rect -30483 7758 -30474 7794
rect -30438 7758 -30429 7794
rect -30483 7749 -30429 7758
rect -30483 7713 -30429 7722
rect -30483 7677 -30474 7713
rect -30438 7677 -30429 7713
rect -30483 7659 -30429 7677
rect -30483 7632 -30429 7641
rect -30483 7596 -30474 7632
rect -30438 7596 -30429 7632
rect -30483 7587 -30429 7596
rect -29673 8163 -29619 8172
rect -29673 8127 -29664 8163
rect -29628 8127 -29619 8163
rect -29673 8118 -29619 8127
rect -29673 8064 -29619 8073
rect -29673 8028 -29664 8064
rect -29628 8028 -29619 8064
rect -29673 8019 -29619 8028
rect -28791 8235 -28737 8244
rect -28791 8199 -28782 8235
rect -28746 8199 -28737 8235
rect -28791 8190 -28737 8199
rect -29673 7992 -29619 8001
rect -29673 7956 -29664 7992
rect -29628 7956 -29619 7992
rect -29673 7947 -29619 7956
rect -29673 7875 -29619 7884
rect -29673 7839 -29664 7875
rect -29628 7839 -29619 7875
rect -29673 7821 -29619 7839
rect -29673 7794 -29619 7803
rect -29673 7758 -29664 7794
rect -29628 7758 -29619 7794
rect -29673 7749 -29619 7758
rect -29673 7713 -29619 7722
rect -29673 7677 -29664 7713
rect -29628 7677 -29619 7713
rect -29673 7659 -29619 7677
rect -29673 7632 -29619 7641
rect -29673 7596 -29664 7632
rect -29628 7596 -29619 7632
rect -29673 7587 -29619 7596
rect -28791 8163 -28737 8172
rect -28791 8127 -28782 8163
rect -28746 8127 -28737 8163
rect -28791 8118 -28737 8127
rect -28791 8064 -28737 8073
rect -28791 8028 -28782 8064
rect -28746 8028 -28737 8064
rect -28791 8019 -28737 8028
rect -28791 7992 -28737 8001
rect -28791 7956 -28782 7992
rect -28746 7956 -28737 7992
rect -28791 7947 -28737 7956
rect -28791 7875 -28737 7884
rect -28791 7839 -28782 7875
rect -28746 7839 -28737 7875
rect -28791 7821 -28737 7839
rect -28791 7794 -28737 7803
rect -28791 7758 -28782 7794
rect -28746 7758 -28737 7794
rect -28791 7749 -28737 7758
rect -28791 7713 -28737 7722
rect -28791 7677 -28782 7713
rect -28746 7677 -28737 7713
rect -28791 7659 -28737 7677
rect -28791 7632 -28737 7641
rect -28791 7596 -28782 7632
rect -28746 7596 -28737 7632
rect -28791 7587 -28737 7596
rect -29916 7146 -29871 7155
rect -29916 7128 -29907 7146
rect -29880 7128 -29871 7146
rect -29853 7128 -29835 7155
rect -29808 7128 -29799 7155
rect -30366 7092 -30330 7101
rect -30366 7074 -30357 7092
rect -30339 7074 -30330 7092
rect -30312 7074 -30168 7101
rect -30150 7083 -30141 7101
rect -30123 7083 -30114 7101
rect -30150 7074 -30114 7083
rect -29340 7155 -29304 7164
rect -29340 7137 -29331 7155
rect -29313 7137 -29304 7155
rect -29286 7137 -29142 7164
rect -29124 7146 -29115 7164
rect -29097 7146 -29088 7164
rect -29124 7137 -29088 7146
rect -28890 7209 -28845 7218
rect -28890 7191 -28881 7209
rect -28854 7191 -28845 7209
rect -28827 7191 -28809 7218
rect -28782 7191 -28773 7218
rect -29691 6732 -29682 6750
rect -29664 6732 -29655 6750
rect -29691 6723 -29655 6732
rect -29637 6732 -29628 6750
rect -29637 6723 -29610 6732
rect -29601 6732 -29592 6750
rect -29574 6732 -29565 6750
rect -29601 6723 -29565 6732
rect -29547 6732 -29538 6750
rect -29547 6723 -29520 6732
rect -29475 6732 -29466 6750
rect -29448 6732 -29439 6750
rect -29475 6723 -29439 6732
rect -29421 6732 -29412 6750
rect -29394 6732 -29385 6750
rect -29421 6723 -29385 6732
rect -30483 6120 -30429 6129
rect -30483 6084 -30474 6120
rect -30438 6084 -30429 6120
rect -30483 6075 -30429 6084
rect -30483 6048 -30429 6057
rect -30483 6012 -30474 6048
rect -30438 6012 -30429 6048
rect -30483 6003 -30429 6012
rect -30483 5949 -30429 5958
rect -30483 5913 -30474 5949
rect -30438 5913 -30429 5949
rect -30483 5904 -30429 5913
rect -29673 6120 -29619 6129
rect -29673 6084 -29664 6120
rect -29628 6084 -29619 6120
rect -29673 6075 -29619 6084
rect -30483 5877 -30429 5886
rect -30483 5841 -30474 5877
rect -30438 5841 -30429 5877
rect -30483 5832 -30429 5841
rect -30483 5760 -30429 5769
rect -30483 5724 -30474 5760
rect -30438 5724 -30429 5760
rect -30483 5706 -30429 5724
rect -30483 5679 -30429 5688
rect -30483 5643 -30474 5679
rect -30438 5643 -30429 5679
rect -30483 5634 -30429 5643
rect -30483 5598 -30429 5607
rect -30483 5562 -30474 5598
rect -30438 5562 -30429 5598
rect -30483 5544 -30429 5562
rect -30483 5517 -30429 5526
rect -30483 5481 -30474 5517
rect -30438 5481 -30429 5517
rect -30483 5472 -30429 5481
rect -29673 6048 -29619 6057
rect -29673 6012 -29664 6048
rect -29628 6012 -29619 6048
rect -29673 6003 -29619 6012
rect -29673 5949 -29619 5958
rect -29673 5913 -29664 5949
rect -29628 5913 -29619 5949
rect -29673 5904 -29619 5913
rect -28791 6120 -28737 6129
rect -28791 6084 -28782 6120
rect -28746 6084 -28737 6120
rect -28791 6075 -28737 6084
rect -29673 5877 -29619 5886
rect -29673 5841 -29664 5877
rect -29628 5841 -29619 5877
rect -29673 5832 -29619 5841
rect -29673 5760 -29619 5769
rect -29673 5724 -29664 5760
rect -29628 5724 -29619 5760
rect -29673 5706 -29619 5724
rect -29673 5679 -29619 5688
rect -29673 5643 -29664 5679
rect -29628 5643 -29619 5679
rect -29673 5634 -29619 5643
rect -29673 5598 -29619 5607
rect -29673 5562 -29664 5598
rect -29628 5562 -29619 5598
rect -29673 5544 -29619 5562
rect -29673 5517 -29619 5526
rect -29673 5481 -29664 5517
rect -29628 5481 -29619 5517
rect -29673 5472 -29619 5481
rect -28791 6048 -28737 6057
rect -28791 6012 -28782 6048
rect -28746 6012 -28737 6048
rect -28791 6003 -28737 6012
rect -28791 5949 -28737 5958
rect -28791 5913 -28782 5949
rect -28746 5913 -28737 5949
rect -28791 5904 -28737 5913
rect -28791 5877 -28737 5886
rect -28791 5841 -28782 5877
rect -28746 5841 -28737 5877
rect -28791 5832 -28737 5841
rect -28791 5760 -28737 5769
rect -28791 5724 -28782 5760
rect -28746 5724 -28737 5760
rect -28791 5706 -28737 5724
rect -28791 5679 -28737 5688
rect -28791 5643 -28782 5679
rect -28746 5643 -28737 5679
rect -28791 5634 -28737 5643
rect -28791 5598 -28737 5607
rect -28791 5562 -28782 5598
rect -28746 5562 -28737 5598
rect -28791 5544 -28737 5562
rect -28791 5517 -28737 5526
rect -28791 5481 -28782 5517
rect -28746 5481 -28737 5517
rect -28791 5472 -28737 5481
rect -29916 5031 -29871 5040
rect -29916 5013 -29907 5031
rect -29880 5013 -29871 5031
rect -29853 5013 -29835 5040
rect -29808 5013 -29799 5040
rect -30366 4977 -30330 4986
rect -30366 4959 -30357 4977
rect -30339 4959 -30330 4977
rect -30312 4959 -30168 4986
rect -30150 4968 -30141 4986
rect -30123 4968 -30114 4986
rect -30150 4959 -30114 4968
rect -29340 5040 -29304 5049
rect -29340 5022 -29331 5040
rect -29313 5022 -29304 5040
rect -29286 5022 -29142 5049
rect -29124 5031 -29115 5049
rect -29097 5031 -29088 5049
rect -29124 5022 -29088 5031
rect -28890 5094 -28845 5103
rect -28890 5076 -28881 5094
rect -28854 5076 -28845 5094
rect -28827 5076 -28809 5103
rect -28782 5076 -28773 5103
rect -29691 4617 -29682 4635
rect -29664 4617 -29655 4635
rect -29691 4608 -29655 4617
rect -29637 4617 -29628 4635
rect -29637 4608 -29610 4617
rect -29601 4617 -29592 4635
rect -29574 4617 -29565 4635
rect -29601 4608 -29565 4617
rect -29547 4617 -29538 4635
rect -29547 4608 -29520 4617
rect -29475 4617 -29466 4635
rect -29448 4617 -29439 4635
rect -29475 4608 -29439 4617
rect -29421 4617 -29412 4635
rect -29394 4617 -29385 4635
rect -29421 4608 -29385 4617
rect -30483 4185 -30429 4194
rect -30483 4149 -30474 4185
rect -30438 4149 -30429 4185
rect -30483 4140 -30429 4149
rect -30483 4113 -30429 4122
rect -30483 4077 -30474 4113
rect -30438 4077 -30429 4113
rect -30483 4068 -30429 4077
rect -30483 4014 -30429 4023
rect -30483 3978 -30474 4014
rect -30438 3978 -30429 4014
rect -30483 3969 -30429 3978
rect -29673 4185 -29619 4194
rect -29673 4149 -29664 4185
rect -29628 4149 -29619 4185
rect -29673 4140 -29619 4149
rect -30483 3942 -30429 3951
rect -30483 3906 -30474 3942
rect -30438 3906 -30429 3942
rect -30483 3897 -30429 3906
rect -30483 3825 -30429 3834
rect -30483 3789 -30474 3825
rect -30438 3789 -30429 3825
rect -30483 3771 -30429 3789
rect -30483 3744 -30429 3753
rect -30483 3708 -30474 3744
rect -30438 3708 -30429 3744
rect -30483 3699 -30429 3708
rect -30483 3663 -30429 3672
rect -30483 3627 -30474 3663
rect -30438 3627 -30429 3663
rect -30483 3609 -30429 3627
rect -30483 3582 -30429 3591
rect -30483 3546 -30474 3582
rect -30438 3546 -30429 3582
rect -30483 3537 -30429 3546
rect -29673 4113 -29619 4122
rect -29673 4077 -29664 4113
rect -29628 4077 -29619 4113
rect -29673 4068 -29619 4077
rect -29673 4014 -29619 4023
rect -29673 3978 -29664 4014
rect -29628 3978 -29619 4014
rect -29673 3969 -29619 3978
rect -28791 4185 -28737 4194
rect -28791 4149 -28782 4185
rect -28746 4149 -28737 4185
rect -28791 4140 -28737 4149
rect -29673 3942 -29619 3951
rect -29673 3906 -29664 3942
rect -29628 3906 -29619 3942
rect -29673 3897 -29619 3906
rect -29673 3825 -29619 3834
rect -29673 3789 -29664 3825
rect -29628 3789 -29619 3825
rect -29673 3771 -29619 3789
rect -29673 3744 -29619 3753
rect -29673 3708 -29664 3744
rect -29628 3708 -29619 3744
rect -29673 3699 -29619 3708
rect -29673 3663 -29619 3672
rect -29673 3627 -29664 3663
rect -29628 3627 -29619 3663
rect -29673 3609 -29619 3627
rect -29673 3582 -29619 3591
rect -29673 3546 -29664 3582
rect -29628 3546 -29619 3582
rect -29673 3537 -29619 3546
rect -28791 4113 -28737 4122
rect -28791 4077 -28782 4113
rect -28746 4077 -28737 4113
rect -28791 4068 -28737 4077
rect -28791 4014 -28737 4023
rect -28791 3978 -28782 4014
rect -28746 3978 -28737 4014
rect -28791 3969 -28737 3978
rect -28791 3942 -28737 3951
rect -28791 3906 -28782 3942
rect -28746 3906 -28737 3942
rect -28791 3897 -28737 3906
rect -28791 3825 -28737 3834
rect -28791 3789 -28782 3825
rect -28746 3789 -28737 3825
rect -28791 3771 -28737 3789
rect -28791 3744 -28737 3753
rect -28791 3708 -28782 3744
rect -28746 3708 -28737 3744
rect -28791 3699 -28737 3708
rect -28791 3663 -28737 3672
rect -28791 3627 -28782 3663
rect -28746 3627 -28737 3663
rect -28791 3609 -28737 3627
rect -28791 3582 -28737 3591
rect -28791 3546 -28782 3582
rect -28746 3546 -28737 3582
rect -28791 3537 -28737 3546
rect -29916 3096 -29871 3105
rect -29916 3078 -29907 3096
rect -29880 3078 -29871 3096
rect -29853 3078 -29835 3105
rect -29808 3078 -29799 3105
rect -30366 3042 -30330 3051
rect -30366 3024 -30357 3042
rect -30339 3024 -30330 3042
rect -30312 3024 -30168 3051
rect -30150 3033 -30141 3051
rect -30123 3033 -30114 3051
rect -30150 3024 -30114 3033
rect -29340 3105 -29304 3114
rect -29340 3087 -29331 3105
rect -29313 3087 -29304 3105
rect -29286 3087 -29142 3114
rect -29124 3096 -29115 3114
rect -29097 3096 -29088 3114
rect -29124 3087 -29088 3096
rect -28890 3159 -28845 3168
rect -28890 3141 -28881 3159
rect -28854 3141 -28845 3159
rect -28827 3141 -28809 3168
rect -28782 3141 -28773 3168
rect -29691 2682 -29682 2700
rect -29664 2682 -29655 2700
rect -29691 2673 -29655 2682
rect -29637 2682 -29628 2700
rect -29637 2673 -29610 2682
rect -29601 2682 -29592 2700
rect -29574 2682 -29565 2700
rect -29601 2673 -29565 2682
rect -29547 2682 -29538 2700
rect -29547 2673 -29520 2682
rect -29475 2682 -29466 2700
rect -29448 2682 -29439 2700
rect -29475 2673 -29439 2682
rect -29421 2682 -29412 2700
rect -29394 2682 -29385 2700
rect -29421 2673 -29385 2682
rect -30123 495 -30069 504
rect -30123 459 -30114 495
rect -30078 459 -30069 495
rect -30123 450 -30069 459
rect -30123 423 -30069 432
rect -30123 387 -30114 423
rect -30078 387 -30069 423
rect -30123 378 -30069 387
rect -30123 324 -30069 333
rect -30123 288 -30114 324
rect -30078 288 -30069 324
rect -30123 279 -30069 288
rect -29520 261 -29475 270
rect -30123 252 -30069 261
rect -30123 216 -30114 252
rect -30078 216 -30069 252
rect -30123 207 -30069 216
rect -29520 243 -29511 261
rect -29484 243 -29475 261
rect -29457 243 -29439 270
rect -29412 243 -29403 270
rect -30123 135 -30069 144
rect -30123 99 -30114 135
rect -30078 99 -30069 135
rect -30123 81 -30069 99
rect -30123 54 -30069 63
rect -30123 18 -30114 54
rect -30078 18 -30069 54
rect -30123 9 -30069 18
rect -30123 -27 -30069 -18
rect -30123 -63 -30114 -27
rect -30078 -63 -30069 -27
rect -30123 -81 -30069 -63
rect -30123 -108 -30069 -99
rect -30123 -144 -30114 -108
rect -30078 -144 -30069 -108
rect -30123 -153 -30069 -144
rect -29151 -45 -29106 -36
rect -29151 -63 -29142 -45
rect -29115 -63 -29106 -45
rect -29088 -63 -29070 -36
rect -29043 -63 -29034 -36
rect -28314 -9 -28269 0
rect -28314 -27 -28305 -9
rect -28278 -27 -28269 -9
rect -28251 -27 -28233 0
rect -28206 -27 -28197 0
rect -28764 -63 -28728 -54
rect -28764 -81 -28755 -63
rect -28737 -81 -28728 -63
rect -28710 -81 -28620 -54
rect -28611 -81 -28566 -54
rect -28548 -72 -28539 -54
rect -28521 -72 -28512 -54
rect -28548 -81 -28512 -72
rect -33444 -423 -33399 -414
rect -33444 -441 -33435 -423
rect -33408 -441 -33399 -423
rect -33381 -441 -33363 -414
rect -33336 -441 -33327 -414
rect -33894 -477 -33858 -468
rect -33894 -495 -33885 -477
rect -33867 -495 -33858 -477
rect -33840 -495 -33696 -468
rect -33678 -486 -33669 -468
rect -33651 -486 -33642 -468
rect -33678 -495 -33642 -486
rect -30123 -450 -30069 -441
rect -30123 -486 -30114 -450
rect -30078 -486 -30069 -450
rect -30123 -495 -30069 -486
rect -33444 -918 -33399 -909
rect -33444 -936 -33435 -918
rect -33408 -936 -33399 -918
rect -33381 -936 -33363 -909
rect -33336 -936 -33327 -909
rect -33894 -972 -33858 -963
rect -33894 -990 -33885 -972
rect -33867 -990 -33858 -972
rect -33840 -990 -33696 -963
rect -33678 -981 -33669 -963
rect -33651 -981 -33642 -963
rect -33678 -990 -33642 -981
rect -34461 -1224 -34452 -1206
rect -34434 -1224 -34425 -1206
rect -34461 -1233 -34425 -1224
rect -34407 -1224 -34398 -1206
rect -34407 -1233 -34380 -1224
rect -34371 -1224 -34362 -1206
rect -34344 -1224 -34335 -1206
rect -34371 -1233 -34335 -1224
rect -34317 -1224 -34308 -1206
rect -34317 -1233 -34290 -1224
rect -34245 -1224 -34236 -1206
rect -34218 -1224 -34209 -1206
rect -34245 -1233 -34209 -1224
rect -34191 -1224 -34182 -1206
rect -34164 -1224 -34155 -1206
rect -34191 -1233 -34155 -1224
rect -33444 -1332 -33399 -1323
rect -33444 -1350 -33435 -1332
rect -33408 -1350 -33399 -1332
rect -33381 -1350 -33363 -1323
rect -33336 -1350 -33327 -1323
rect -33894 -1386 -33858 -1377
rect -33894 -1404 -33885 -1386
rect -33867 -1404 -33858 -1386
rect -33840 -1404 -33696 -1377
rect -33678 -1395 -33669 -1377
rect -33651 -1395 -33642 -1377
rect -33678 -1404 -33642 -1395
rect -33444 -1863 -33399 -1854
rect -33444 -1881 -33435 -1863
rect -33408 -1881 -33399 -1863
rect -33381 -1881 -33363 -1854
rect -33336 -1881 -33327 -1854
rect -33894 -1917 -33858 -1908
rect -33894 -1935 -33885 -1917
rect -33867 -1935 -33858 -1917
rect -33840 -1935 -33696 -1908
rect -33678 -1926 -33669 -1908
rect -33651 -1926 -33642 -1908
rect -33678 -1935 -33642 -1926
rect -33444 -2430 -33399 -2421
rect -33444 -2448 -33435 -2430
rect -33408 -2448 -33399 -2430
rect -33381 -2448 -33363 -2421
rect -33336 -2448 -33327 -2421
rect -33894 -2484 -33858 -2475
rect -33894 -2502 -33885 -2484
rect -33867 -2502 -33858 -2484
rect -33840 -2502 -33696 -2475
rect -33678 -2493 -33669 -2475
rect -33651 -2493 -33642 -2475
rect -33678 -2502 -33642 -2493
rect -33444 -2925 -33399 -2916
rect -33444 -2943 -33435 -2925
rect -33408 -2943 -33399 -2925
rect -33381 -2943 -33363 -2916
rect -33336 -2943 -33327 -2916
rect -33894 -2979 -33858 -2970
rect -33894 -2997 -33885 -2979
rect -33867 -2997 -33858 -2979
rect -33840 -2997 -33696 -2970
rect -33678 -2988 -33669 -2970
rect -33651 -2988 -33642 -2970
rect -33678 -2997 -33642 -2988
rect -33444 -3339 -33399 -3330
rect -33444 -3357 -33435 -3339
rect -33408 -3357 -33399 -3339
rect -33381 -3357 -33363 -3330
rect -33336 -3357 -33327 -3330
rect -33894 -3393 -33858 -3384
rect -33894 -3411 -33885 -3393
rect -33867 -3411 -33858 -3393
rect -33840 -3411 -33696 -3384
rect -33678 -3402 -33669 -3384
rect -33651 -3402 -33642 -3384
rect -33678 -3411 -33642 -3402
rect -33444 -3870 -33399 -3861
rect -33444 -3888 -33435 -3870
rect -33408 -3888 -33399 -3870
rect -33381 -3888 -33363 -3861
rect -33336 -3888 -33327 -3861
rect -33894 -3924 -33858 -3915
rect -33894 -3942 -33885 -3924
rect -33867 -3942 -33858 -3924
rect -33840 -3942 -33696 -3915
rect -33678 -3933 -33669 -3915
rect -33651 -3933 -33642 -3915
rect -33678 -3942 -33642 -3933
rect -30123 -522 -30069 -513
rect -30123 -558 -30114 -522
rect -30078 -558 -30069 -522
rect -30123 -567 -30069 -558
rect -30123 -621 -30069 -612
rect -30123 -657 -30114 -621
rect -30078 -657 -30069 -621
rect -30123 -666 -30069 -657
rect -29520 -684 -29475 -675
rect -30123 -693 -30069 -684
rect -30123 -729 -30114 -693
rect -30078 -729 -30069 -693
rect -30123 -738 -30069 -729
rect -29520 -702 -29511 -684
rect -29484 -702 -29475 -684
rect -29457 -702 -29439 -675
rect -29412 -702 -29403 -675
rect -30123 -810 -30069 -801
rect -30123 -846 -30114 -810
rect -30078 -846 -30069 -810
rect -30123 -864 -30069 -846
rect -30123 -891 -30069 -882
rect -30123 -927 -30114 -891
rect -30078 -927 -30069 -891
rect -30123 -936 -30069 -927
rect -29169 -855 -29124 -846
rect -29169 -873 -29160 -855
rect -29133 -873 -29124 -855
rect -29106 -873 -29088 -846
rect -29061 -873 -29052 -846
rect -28386 -819 -28341 -810
rect -28386 -837 -28377 -819
rect -28350 -837 -28341 -819
rect -28323 -837 -28305 -810
rect -28278 -837 -28269 -810
rect -27558 -819 -27513 -810
rect -27558 -837 -27549 -819
rect -27522 -837 -27513 -819
rect -27495 -837 -27477 -810
rect -27450 -837 -27441 -810
rect -28836 -873 -28800 -864
rect -28836 -891 -28827 -873
rect -28809 -891 -28800 -873
rect -28782 -891 -28692 -864
rect -28683 -891 -28638 -864
rect -28620 -882 -28611 -864
rect -28593 -882 -28584 -864
rect -28620 -891 -28584 -882
rect -28008 -873 -27972 -864
rect -28008 -891 -27999 -873
rect -27981 -891 -27972 -873
rect -27954 -891 -27810 -864
rect -27792 -882 -27783 -864
rect -27765 -882 -27756 -864
rect -27792 -891 -27756 -882
rect -27135 -882 -27126 -864
rect -27108 -882 -27090 -864
rect -27135 -891 -27090 -882
rect -27072 -882 -27063 -864
rect -27072 -891 -27045 -882
rect -27036 -882 -27027 -864
rect -27009 -882 -27000 -864
rect -27036 -891 -27000 -882
rect -26982 -882 -26973 -864
rect -26982 -891 -26955 -882
rect -26946 -882 -26937 -864
rect -26919 -882 -26910 -864
rect -26946 -891 -26910 -882
rect -26892 -882 -26883 -864
rect -26892 -891 -26865 -882
rect -26856 -882 -26847 -864
rect -26829 -882 -26820 -864
rect -26856 -891 -26820 -882
rect -26802 -882 -26793 -864
rect -26802 -891 -26775 -882
rect -26730 -882 -26721 -864
rect -26703 -882 -26694 -864
rect -26730 -891 -26694 -882
rect -26676 -882 -26667 -864
rect -26649 -882 -26640 -864
rect -26676 -891 -26640 -882
rect -30123 -972 -30069 -963
rect -30123 -1008 -30114 -972
rect -30078 -1008 -30069 -972
rect -30123 -1026 -30069 -1008
rect -30123 -1053 -30069 -1044
rect -30123 -1089 -30114 -1053
rect -30078 -1089 -30069 -1053
rect -30123 -1098 -30069 -1089
rect -30123 -1467 -30069 -1458
rect -30123 -1503 -30114 -1467
rect -30078 -1503 -30069 -1467
rect -30123 -1512 -30069 -1503
rect -30123 -1539 -30069 -1530
rect -30123 -1575 -30114 -1539
rect -30078 -1575 -30069 -1539
rect -30123 -1584 -30069 -1575
rect -30123 -1638 -30069 -1629
rect -30123 -1674 -30114 -1638
rect -30078 -1674 -30069 -1638
rect -30123 -1683 -30069 -1674
rect -29520 -1701 -29475 -1692
rect -30123 -1710 -30069 -1701
rect -30123 -1746 -30114 -1710
rect -30078 -1746 -30069 -1710
rect -30123 -1755 -30069 -1746
rect -29520 -1719 -29511 -1701
rect -29484 -1719 -29475 -1701
rect -29457 -1719 -29439 -1692
rect -29412 -1719 -29403 -1692
rect -29187 -1701 -29142 -1692
rect -29187 -1719 -29178 -1701
rect -29151 -1719 -29142 -1701
rect -29124 -1719 -29106 -1692
rect -29079 -1719 -29070 -1692
rect -28683 -1701 -28674 -1674
rect -28647 -1701 -28638 -1674
rect -28620 -1701 -28512 -1674
rect -28494 -1701 -28368 -1674
rect -28350 -1701 -28242 -1674
rect -28224 -1701 -28107 -1674
rect -28089 -1701 -28053 -1674
rect -28026 -1701 -27954 -1674
rect -27900 -1701 -27882 -1674
rect -27855 -1701 -27846 -1674
rect -27828 -1701 -27819 -1674
rect -27792 -1701 -27783 -1674
rect -30123 -1827 -30069 -1818
rect -30123 -1863 -30114 -1827
rect -30078 -1863 -30069 -1827
rect -30123 -1881 -30069 -1863
rect -30123 -1908 -30069 -1899
rect -30123 -1944 -30114 -1908
rect -30078 -1944 -30069 -1908
rect -30123 -1953 -30069 -1944
rect -30123 -1989 -30069 -1980
rect -30123 -2025 -30114 -1989
rect -30078 -2025 -30069 -1989
rect -30123 -2043 -30069 -2025
rect -30123 -2070 -30069 -2061
rect -30123 -2106 -30114 -2070
rect -30078 -2106 -30069 -2070
rect -30123 -2115 -30069 -2106
rect -30123 -2763 -30069 -2754
rect -30123 -2799 -30114 -2763
rect -30078 -2799 -30069 -2763
rect -30123 -2808 -30069 -2799
rect -30123 -2835 -30069 -2826
rect -30123 -2871 -30114 -2835
rect -30078 -2871 -30069 -2835
rect -30123 -2880 -30069 -2871
rect -30123 -2934 -30069 -2925
rect -30123 -2970 -30114 -2934
rect -30078 -2970 -30069 -2934
rect -30123 -2979 -30069 -2970
rect -29520 -2997 -29475 -2988
rect -30123 -3006 -30069 -2997
rect -30123 -3042 -30114 -3006
rect -30078 -3042 -30069 -3006
rect -30123 -3051 -30069 -3042
rect -29520 -3015 -29511 -2997
rect -29484 -3015 -29475 -2997
rect -29457 -3015 -29439 -2988
rect -29412 -3015 -29403 -2988
rect -29241 -2997 -29196 -2988
rect -29241 -3015 -29232 -2997
rect -29205 -3015 -29196 -2997
rect -29178 -3015 -29160 -2988
rect -29133 -3015 -29124 -2988
rect -28836 -2997 -28827 -2970
rect -28800 -2997 -28791 -2970
rect -28773 -2997 -28665 -2970
rect -28647 -2997 -28521 -2970
rect -28503 -2997 -28395 -2970
rect -28377 -2997 -28260 -2970
rect -28242 -2997 -28206 -2970
rect -28179 -2997 -28107 -2970
rect -28053 -2997 -28035 -2970
rect -28008 -2997 -27999 -2970
rect -27981 -2997 -27972 -2970
rect -27945 -2997 -27936 -2970
rect -30123 -3123 -30069 -3114
rect -30123 -3159 -30114 -3123
rect -30078 -3159 -30069 -3123
rect -30123 -3177 -30069 -3159
rect -30123 -3204 -30069 -3195
rect -30123 -3240 -30114 -3204
rect -30078 -3240 -30069 -3204
rect -30123 -3249 -30069 -3240
rect -30123 -3285 -30069 -3276
rect -30123 -3321 -30114 -3285
rect -30078 -3321 -30069 -3285
rect -30123 -3339 -30069 -3321
rect -30123 -3366 -30069 -3357
rect -30123 -3402 -30114 -3366
rect -30078 -3402 -30069 -3366
rect -30123 -3411 -30069 -3402
rect -30123 -3834 -30069 -3825
rect -30123 -3870 -30114 -3834
rect -30078 -3870 -30069 -3834
rect -30123 -3879 -30069 -3870
rect -30123 -3906 -30069 -3897
rect -30123 -3942 -30114 -3906
rect -30078 -3942 -30069 -3906
rect -30123 -3951 -30069 -3942
rect -30123 -4005 -30069 -3996
rect -30123 -4041 -30114 -4005
rect -30078 -4041 -30069 -4005
rect -30123 -4050 -30069 -4041
rect -29520 -4068 -29475 -4059
rect -30123 -4077 -30069 -4068
rect -30123 -4113 -30114 -4077
rect -30078 -4113 -30069 -4077
rect -30123 -4122 -30069 -4113
rect -29520 -4086 -29511 -4068
rect -29484 -4086 -29475 -4068
rect -29457 -4086 -29439 -4059
rect -29412 -4086 -29403 -4059
rect -30123 -4194 -30069 -4185
rect -30123 -4230 -30114 -4194
rect -30078 -4230 -30069 -4194
rect -30123 -4248 -30069 -4230
rect -30123 -4275 -30069 -4266
rect -30123 -4311 -30114 -4275
rect -30078 -4311 -30069 -4275
rect -30123 -4320 -30069 -4311
rect -30123 -4356 -30069 -4347
rect -30123 -4392 -30114 -4356
rect -30078 -4392 -30069 -4356
rect -30123 -4410 -30069 -4392
rect -30123 -4437 -30069 -4428
rect -30123 -4473 -30114 -4437
rect -30078 -4473 -30069 -4437
rect -30123 -4482 -30069 -4473
rect -29151 -4374 -29106 -4365
rect -29151 -4392 -29142 -4374
rect -29115 -4392 -29106 -4374
rect -29088 -4392 -29070 -4365
rect -29043 -4392 -29034 -4365
rect -28314 -4338 -28269 -4329
rect -28314 -4356 -28305 -4338
rect -28278 -4356 -28269 -4338
rect -28251 -4356 -28233 -4329
rect -28206 -4356 -28197 -4329
rect -28764 -4392 -28728 -4383
rect -28764 -4410 -28755 -4392
rect -28737 -4410 -28728 -4392
rect -28710 -4410 -28620 -4383
rect -28611 -4410 -28566 -4383
rect -28548 -4401 -28539 -4383
rect -28521 -4401 -28512 -4383
rect -28548 -4410 -28512 -4401
rect -30123 -4779 -30069 -4770
rect -30123 -4815 -30114 -4779
rect -30078 -4815 -30069 -4779
rect -30123 -4824 -30069 -4815
rect -30123 -4851 -30069 -4842
rect -30123 -4887 -30114 -4851
rect -30078 -4887 -30069 -4851
rect -30123 -4896 -30069 -4887
rect -30123 -4950 -30069 -4941
rect -30123 -4986 -30114 -4950
rect -30078 -4986 -30069 -4950
rect -30123 -4995 -30069 -4986
rect -29520 -5013 -29475 -5004
rect -30123 -5022 -30069 -5013
rect -30123 -5058 -30114 -5022
rect -30078 -5058 -30069 -5022
rect -30123 -5067 -30069 -5058
rect -29520 -5031 -29511 -5013
rect -29484 -5031 -29475 -5013
rect -29457 -5031 -29439 -5004
rect -29412 -5031 -29403 -5004
rect -30123 -5139 -30069 -5130
rect -30123 -5175 -30114 -5139
rect -30078 -5175 -30069 -5139
rect -30123 -5193 -30069 -5175
rect -30123 -5220 -30069 -5211
rect -30123 -5256 -30114 -5220
rect -30078 -5256 -30069 -5220
rect -30123 -5265 -30069 -5256
rect -29169 -5184 -29124 -5175
rect -29169 -5202 -29160 -5184
rect -29133 -5202 -29124 -5184
rect -29106 -5202 -29088 -5175
rect -29061 -5202 -29052 -5175
rect -28386 -5148 -28341 -5139
rect -28386 -5166 -28377 -5148
rect -28350 -5166 -28341 -5148
rect -28323 -5166 -28305 -5139
rect -28278 -5166 -28269 -5139
rect -27558 -5148 -27513 -5139
rect -27558 -5166 -27549 -5148
rect -27522 -5166 -27513 -5148
rect -27495 -5166 -27477 -5139
rect -27450 -5166 -27441 -5139
rect -28836 -5202 -28800 -5193
rect -28836 -5220 -28827 -5202
rect -28809 -5220 -28800 -5202
rect -28782 -5220 -28692 -5193
rect -28683 -5220 -28638 -5193
rect -28620 -5211 -28611 -5193
rect -28593 -5211 -28584 -5193
rect -28620 -5220 -28584 -5211
rect -28008 -5202 -27972 -5193
rect -28008 -5220 -27999 -5202
rect -27981 -5220 -27972 -5202
rect -27954 -5220 -27810 -5193
rect -27792 -5211 -27783 -5193
rect -27765 -5211 -27756 -5193
rect -27792 -5220 -27756 -5211
rect -27135 -5211 -27126 -5193
rect -27108 -5211 -27090 -5193
rect -27135 -5220 -27090 -5211
rect -27072 -5211 -27063 -5193
rect -27072 -5220 -27045 -5211
rect -27036 -5211 -27027 -5193
rect -27009 -5211 -27000 -5193
rect -27036 -5220 -27000 -5211
rect -26982 -5211 -26973 -5193
rect -26982 -5220 -26955 -5211
rect -26946 -5211 -26937 -5193
rect -26919 -5211 -26910 -5193
rect -26946 -5220 -26910 -5211
rect -26892 -5211 -26883 -5193
rect -26892 -5220 -26865 -5211
rect -26856 -5211 -26847 -5193
rect -26829 -5211 -26820 -5193
rect -26856 -5220 -26820 -5211
rect -26802 -5211 -26793 -5193
rect -26802 -5220 -26775 -5211
rect -26730 -5211 -26721 -5193
rect -26703 -5211 -26694 -5193
rect -26730 -5220 -26694 -5211
rect -26676 -5211 -26667 -5193
rect -26649 -5211 -26640 -5193
rect -26676 -5220 -26640 -5211
rect -30123 -5301 -30069 -5292
rect -30123 -5337 -30114 -5301
rect -30078 -5337 -30069 -5301
rect -30123 -5355 -30069 -5337
rect -30123 -5382 -30069 -5373
rect -30123 -5418 -30114 -5382
rect -30078 -5418 -30069 -5382
rect -30123 -5427 -30069 -5418
rect -30123 -5796 -30069 -5787
rect -30123 -5832 -30114 -5796
rect -30078 -5832 -30069 -5796
rect -30123 -5841 -30069 -5832
rect -30123 -5868 -30069 -5859
rect -30123 -5904 -30114 -5868
rect -30078 -5904 -30069 -5868
rect -30123 -5913 -30069 -5904
rect -30123 -5967 -30069 -5958
rect -30123 -6003 -30114 -5967
rect -30078 -6003 -30069 -5967
rect -30123 -6012 -30069 -6003
rect -29520 -6030 -29475 -6021
rect -30123 -6039 -30069 -6030
rect -30123 -6075 -30114 -6039
rect -30078 -6075 -30069 -6039
rect -30123 -6084 -30069 -6075
rect -29520 -6048 -29511 -6030
rect -29484 -6048 -29475 -6030
rect -29457 -6048 -29439 -6021
rect -29412 -6048 -29403 -6021
rect -29187 -6030 -29142 -6021
rect -29187 -6048 -29178 -6030
rect -29151 -6048 -29142 -6030
rect -29124 -6048 -29106 -6021
rect -29079 -6048 -29070 -6021
rect -28683 -6030 -28674 -6003
rect -28647 -6030 -28638 -6003
rect -28620 -6030 -28512 -6003
rect -28494 -6030 -28368 -6003
rect -28350 -6030 -28242 -6003
rect -28224 -6030 -28107 -6003
rect -28089 -6030 -28053 -6003
rect -28026 -6030 -27954 -6003
rect -27900 -6030 -27882 -6003
rect -27855 -6030 -27846 -6003
rect -27828 -6030 -27819 -6003
rect -27792 -6030 -27783 -6003
rect -30123 -6156 -30069 -6147
rect -30123 -6192 -30114 -6156
rect -30078 -6192 -30069 -6156
rect -30123 -6210 -30069 -6192
rect -30123 -6237 -30069 -6228
rect -30123 -6273 -30114 -6237
rect -30078 -6273 -30069 -6237
rect -30123 -6282 -30069 -6273
rect -30123 -6318 -30069 -6309
rect -30123 -6354 -30114 -6318
rect -30078 -6354 -30069 -6318
rect -30123 -6372 -30069 -6354
rect -30123 -6399 -30069 -6390
rect -30123 -6435 -30114 -6399
rect -30078 -6435 -30069 -6399
rect -30123 -6444 -30069 -6435
rect -33426 -8280 -33381 -8271
rect -33426 -8298 -33417 -8280
rect -33390 -8298 -33381 -8280
rect -33363 -8298 -33345 -8271
rect -33318 -8298 -33309 -8271
rect -33876 -8334 -33840 -8325
rect -33876 -8352 -33867 -8334
rect -33849 -8352 -33840 -8334
rect -33822 -8352 -33678 -8325
rect -33660 -8343 -33651 -8325
rect -33633 -8343 -33624 -8325
rect -33660 -8352 -33624 -8343
rect -33426 -8775 -33381 -8766
rect -33426 -8793 -33417 -8775
rect -33390 -8793 -33381 -8775
rect -33363 -8793 -33345 -8766
rect -33318 -8793 -33309 -8766
rect -33876 -8829 -33840 -8820
rect -33876 -8847 -33867 -8829
rect -33849 -8847 -33840 -8829
rect -33822 -8847 -33678 -8820
rect -33660 -8838 -33651 -8820
rect -33633 -8838 -33624 -8820
rect -33660 -8847 -33624 -8838
rect -33426 -9189 -33381 -9180
rect -33426 -9207 -33417 -9189
rect -33390 -9207 -33381 -9189
rect -33363 -9207 -33345 -9180
rect -33318 -9207 -33309 -9180
rect -33876 -9243 -33840 -9234
rect -33876 -9261 -33867 -9243
rect -33849 -9261 -33840 -9243
rect -33822 -9261 -33678 -9234
rect -33660 -9252 -33651 -9234
rect -33633 -9252 -33624 -9234
rect -33660 -9261 -33624 -9252
rect -33426 -9720 -33381 -9711
rect -33426 -9738 -33417 -9720
rect -33390 -9738 -33381 -9720
rect -33363 -9738 -33345 -9711
rect -33318 -9738 -33309 -9711
rect -33876 -9774 -33840 -9765
rect -33876 -9792 -33867 -9774
rect -33849 -9792 -33840 -9774
rect -33822 -9792 -33678 -9765
rect -33660 -9783 -33651 -9765
rect -33633 -9783 -33624 -9765
rect -33660 -9792 -33624 -9783
rect -33426 -10197 -33381 -10188
rect -33426 -10215 -33417 -10197
rect -33390 -10215 -33381 -10197
rect -33363 -10215 -33345 -10188
rect -33318 -10215 -33309 -10188
rect -33876 -10251 -33840 -10242
rect -33876 -10269 -33867 -10251
rect -33849 -10269 -33840 -10251
rect -33822 -10269 -33678 -10242
rect -33660 -10260 -33651 -10242
rect -33633 -10260 -33624 -10242
rect -33660 -10269 -33624 -10260
rect -35424 -11619 -35379 -11610
rect -35424 -11637 -35415 -11619
rect -35388 -11637 -35379 -11619
rect -35361 -11637 -35343 -11610
rect -35316 -11637 -35307 -11610
rect -35874 -11673 -35838 -11664
rect -35874 -11691 -35865 -11673
rect -35847 -11691 -35838 -11673
rect -35820 -11691 -35676 -11664
rect -35658 -11682 -35649 -11664
rect -35631 -11682 -35622 -11664
rect -35658 -11691 -35622 -11682
rect -33426 -10692 -33381 -10683
rect -33426 -10710 -33417 -10692
rect -33390 -10710 -33381 -10692
rect -33363 -10710 -33345 -10683
rect -33318 -10710 -33309 -10683
rect -33876 -10746 -33840 -10737
rect -33876 -10764 -33867 -10746
rect -33849 -10764 -33840 -10746
rect -33822 -10764 -33678 -10737
rect -33660 -10755 -33651 -10737
rect -33633 -10755 -33624 -10737
rect -33660 -10764 -33624 -10755
rect -33426 -11106 -33381 -11097
rect -33426 -11124 -33417 -11106
rect -33390 -11124 -33381 -11106
rect -33363 -11124 -33345 -11097
rect -33318 -11124 -33309 -11097
rect -33876 -11160 -33840 -11151
rect -33876 -11178 -33867 -11160
rect -33849 -11178 -33840 -11160
rect -33822 -11178 -33678 -11151
rect -33660 -11169 -33651 -11151
rect -33633 -11169 -33624 -11151
rect -33660 -11178 -33624 -11169
rect -30123 -7092 -30069 -7083
rect -30123 -7128 -30114 -7092
rect -30078 -7128 -30069 -7092
rect -30123 -7137 -30069 -7128
rect -30123 -7164 -30069 -7155
rect -30123 -7200 -30114 -7164
rect -30078 -7200 -30069 -7164
rect -30123 -7209 -30069 -7200
rect -30123 -7263 -30069 -7254
rect -30123 -7299 -30114 -7263
rect -30078 -7299 -30069 -7263
rect -30123 -7308 -30069 -7299
rect -29520 -7326 -29475 -7317
rect -30123 -7335 -30069 -7326
rect -30123 -7371 -30114 -7335
rect -30078 -7371 -30069 -7335
rect -30123 -7380 -30069 -7371
rect -29520 -7344 -29511 -7326
rect -29484 -7344 -29475 -7326
rect -29457 -7344 -29439 -7317
rect -29412 -7344 -29403 -7317
rect -30123 -7452 -30069 -7443
rect -30123 -7488 -30114 -7452
rect -30078 -7488 -30069 -7452
rect -30123 -7506 -30069 -7488
rect -30123 -7533 -30069 -7524
rect -30123 -7569 -30114 -7533
rect -30078 -7569 -30069 -7533
rect -30123 -7578 -30069 -7569
rect -30123 -7614 -30069 -7605
rect -30123 -7650 -30114 -7614
rect -30078 -7650 -30069 -7614
rect -30123 -7668 -30069 -7650
rect -30123 -7695 -30069 -7686
rect -30123 -7731 -30114 -7695
rect -30078 -7731 -30069 -7695
rect -30123 -7740 -30069 -7731
rect -30123 -8631 -30069 -8622
rect -30123 -8667 -30114 -8631
rect -30078 -8667 -30069 -8631
rect -30123 -8676 -30069 -8667
rect -30123 -8703 -30069 -8694
rect -30123 -8739 -30114 -8703
rect -30078 -8739 -30069 -8703
rect -30123 -8748 -30069 -8739
rect -30123 -8802 -30069 -8793
rect -30123 -8838 -30114 -8802
rect -30078 -8838 -30069 -8802
rect -30123 -8847 -30069 -8838
rect -29241 -7326 -29196 -7317
rect -29241 -7344 -29232 -7326
rect -29205 -7344 -29196 -7326
rect -29178 -7344 -29160 -7317
rect -29133 -7344 -29124 -7317
rect -28836 -7326 -28827 -7299
rect -28800 -7326 -28791 -7299
rect -28773 -7326 -28665 -7299
rect -28647 -7326 -28521 -7299
rect -28503 -7326 -28395 -7299
rect -28377 -7326 -28260 -7299
rect -28242 -7326 -28206 -7299
rect -28179 -7326 -28107 -7299
rect -28053 -7326 -28035 -7299
rect -28008 -7326 -27999 -7299
rect -27981 -7326 -27972 -7299
rect -27945 -7326 -27936 -7299
rect -29520 -8865 -29475 -8856
rect -30123 -8874 -30069 -8865
rect -30123 -8910 -30114 -8874
rect -30078 -8910 -30069 -8874
rect -30123 -8919 -30069 -8910
rect -29520 -8883 -29511 -8865
rect -29484 -8883 -29475 -8865
rect -29457 -8883 -29439 -8856
rect -29412 -8883 -29403 -8856
rect -30123 -8991 -30069 -8982
rect -30123 -9027 -30114 -8991
rect -30078 -9027 -30069 -8991
rect -30123 -9045 -30069 -9027
rect -30123 -9072 -30069 -9063
rect -30123 -9108 -30114 -9072
rect -30078 -9108 -30069 -9072
rect -30123 -9117 -30069 -9108
rect -30123 -9153 -30069 -9144
rect -30123 -9189 -30114 -9153
rect -30078 -9189 -30069 -9153
rect -30123 -9207 -30069 -9189
rect -30123 -9234 -30069 -9225
rect -30123 -9270 -30114 -9234
rect -30078 -9270 -30069 -9234
rect -30123 -9279 -30069 -9270
rect -30123 -9576 -30069 -9567
rect -30123 -9612 -30114 -9576
rect -30078 -9612 -30069 -9576
rect -30123 -9621 -30069 -9612
rect -30123 -9648 -30069 -9639
rect -30123 -9684 -30114 -9648
rect -30078 -9684 -30069 -9648
rect -30123 -9693 -30069 -9684
rect -30123 -9747 -30069 -9738
rect -30123 -9783 -30114 -9747
rect -30078 -9783 -30069 -9747
rect -30123 -9792 -30069 -9783
rect -29520 -9810 -29475 -9801
rect -30123 -9819 -30069 -9810
rect -30123 -9855 -30114 -9819
rect -30078 -9855 -30069 -9819
rect -30123 -9864 -30069 -9855
rect -29520 -9828 -29511 -9810
rect -29484 -9828 -29475 -9810
rect -29457 -9828 -29439 -9801
rect -29412 -9828 -29403 -9801
rect -30123 -9936 -30069 -9927
rect -30123 -9972 -30114 -9936
rect -30078 -9972 -30069 -9936
rect -30123 -9990 -30069 -9972
rect -30123 -10017 -30069 -10008
rect -30123 -10053 -30114 -10017
rect -30078 -10053 -30069 -10017
rect -30123 -10062 -30069 -10053
rect -30123 -10098 -30069 -10089
rect -30123 -10134 -30114 -10098
rect -30078 -10134 -30069 -10098
rect -30123 -10152 -30069 -10134
rect -26415 -9873 -26370 -9864
rect -26415 -9891 -26406 -9873
rect -26379 -9891 -26370 -9873
rect -26352 -9891 -26334 -9864
rect -26307 -9891 -26298 -9864
rect -26865 -9927 -26829 -9918
rect -26865 -9945 -26856 -9927
rect -26838 -9945 -26829 -9927
rect -26811 -9945 -26667 -9918
rect -26649 -9936 -26640 -9918
rect -26622 -9936 -26613 -9918
rect -26649 -9945 -26613 -9936
rect -28215 -9981 -28206 -9954
rect -28179 -9981 -28170 -9954
rect -28152 -9981 -28044 -9954
rect -28026 -9981 -27900 -9954
rect -27882 -9981 -27774 -9954
rect -27756 -9981 -27639 -9954
rect -27621 -9981 -27585 -9954
rect -27558 -9981 -27486 -9954
rect -27432 -9981 -27414 -9954
rect -27387 -9981 -27378 -9954
rect -27360 -9981 -27351 -9954
rect -27324 -9981 -27315 -9954
rect -30123 -10179 -30069 -10170
rect -30123 -10215 -30114 -10179
rect -30078 -10215 -30069 -10179
rect -30123 -10224 -30069 -10215
rect -30123 -10593 -30069 -10584
rect -30123 -10629 -30114 -10593
rect -30078 -10629 -30069 -10593
rect -30123 -10638 -30069 -10629
rect -30123 -10665 -30069 -10656
rect -30123 -10701 -30114 -10665
rect -30078 -10701 -30069 -10665
rect -30123 -10710 -30069 -10701
rect -30123 -10764 -30069 -10755
rect -30123 -10800 -30114 -10764
rect -30078 -10800 -30069 -10764
rect -30123 -10809 -30069 -10800
rect -29520 -10827 -29475 -10818
rect -30123 -10836 -30069 -10827
rect -30123 -10872 -30114 -10836
rect -30078 -10872 -30069 -10836
rect -30123 -10881 -30069 -10872
rect -29520 -10845 -29511 -10827
rect -29484 -10845 -29475 -10827
rect -29457 -10845 -29439 -10818
rect -29412 -10845 -29403 -10818
rect -30123 -10953 -30069 -10944
rect -30123 -10989 -30114 -10953
rect -30078 -10989 -30069 -10953
rect -30123 -11007 -30069 -10989
rect -30123 -11034 -30069 -11025
rect -30123 -11070 -30114 -11034
rect -30078 -11070 -30069 -11034
rect -30123 -11079 -30069 -11070
rect -30123 -11115 -30069 -11106
rect -30123 -11151 -30114 -11115
rect -30078 -11151 -30069 -11115
rect -30123 -11169 -30069 -11151
rect -30123 -11196 -30069 -11187
rect -30123 -11232 -30114 -11196
rect -30078 -11232 -30069 -11196
rect -30123 -11241 -30069 -11232
rect -35424 -12087 -35379 -12078
rect -35424 -12105 -35415 -12087
rect -35388 -12105 -35379 -12087
rect -35361 -12105 -35343 -12078
rect -35316 -12105 -35307 -12078
rect -35874 -12141 -35838 -12132
rect -35874 -12159 -35865 -12141
rect -35847 -12159 -35838 -12141
rect -35820 -12159 -35676 -12132
rect -35658 -12150 -35649 -12132
rect -35631 -12150 -35622 -12132
rect -35658 -12159 -35622 -12150
rect -36216 -12276 -36171 -12267
rect -36216 -12294 -36207 -12276
rect -36180 -12294 -36171 -12276
rect -36153 -12294 -36135 -12267
rect -36108 -12294 -36099 -12267
rect -33426 -11637 -33381 -11628
rect -33426 -11655 -33417 -11637
rect -33390 -11655 -33381 -11637
rect -33363 -11655 -33345 -11628
rect -33318 -11655 -33309 -11628
rect -33876 -11691 -33840 -11682
rect -33876 -11709 -33867 -11691
rect -33849 -11709 -33840 -11691
rect -33822 -11709 -33678 -11682
rect -33660 -11700 -33651 -11682
rect -33633 -11700 -33624 -11682
rect -33660 -11709 -33624 -11700
rect -30123 -11889 -30069 -11880
rect -30123 -11925 -30114 -11889
rect -30078 -11925 -30069 -11889
rect -30123 -11934 -30069 -11925
rect -35424 -12528 -35379 -12519
rect -35424 -12546 -35415 -12528
rect -35388 -12546 -35379 -12528
rect -35361 -12546 -35343 -12519
rect -35316 -12546 -35307 -12519
rect -35874 -12582 -35838 -12573
rect -36207 -12600 -36162 -12591
rect -36207 -12618 -36198 -12600
rect -36171 -12618 -36162 -12600
rect -36144 -12618 -36126 -12591
rect -36099 -12618 -36090 -12591
rect -35874 -12600 -35865 -12582
rect -35847 -12600 -35838 -12582
rect -35820 -12600 -35703 -12573
rect -35685 -12600 -35676 -12573
rect -35658 -12591 -35649 -12573
rect -35631 -12591 -35622 -12573
rect -35658 -12600 -35622 -12591
rect -33426 -12501 -33381 -12492
rect -33426 -12519 -33417 -12501
rect -33390 -12519 -33381 -12501
rect -33363 -12519 -33345 -12492
rect -33318 -12519 -33309 -12492
rect -33876 -12555 -33840 -12546
rect -33876 -12573 -33867 -12555
rect -33849 -12573 -33840 -12555
rect -33822 -12573 -33678 -12546
rect -33660 -12564 -33651 -12546
rect -33633 -12564 -33624 -12546
rect -33660 -12573 -33624 -12564
rect -30123 -11961 -30069 -11952
rect -30123 -11997 -30114 -11961
rect -30078 -11997 -30069 -11961
rect -30123 -12006 -30069 -11997
rect -30123 -12060 -30069 -12051
rect -30123 -12096 -30114 -12060
rect -30078 -12096 -30069 -12060
rect -30123 -12105 -30069 -12096
rect -29520 -12123 -29475 -12114
rect -30123 -12132 -30069 -12123
rect -30123 -12168 -30114 -12132
rect -30078 -12168 -30069 -12132
rect -30123 -12177 -30069 -12168
rect -29520 -12141 -29511 -12123
rect -29484 -12141 -29475 -12123
rect -29457 -12141 -29439 -12114
rect -29412 -12141 -29403 -12114
rect -30123 -12249 -30069 -12240
rect -30123 -12285 -30114 -12249
rect -30078 -12285 -30069 -12249
rect -30123 -12303 -30069 -12285
rect -30123 -12330 -30069 -12321
rect -30123 -12366 -30114 -12330
rect -30078 -12366 -30069 -12330
rect -30123 -12375 -30069 -12366
rect -30123 -12411 -30069 -12402
rect -30123 -12447 -30114 -12411
rect -30078 -12447 -30069 -12411
rect -30123 -12465 -30069 -12447
rect -30123 -12492 -30069 -12483
rect -30123 -12528 -30114 -12492
rect -30078 -12528 -30069 -12492
rect -30123 -12537 -30069 -12528
rect -35424 -12942 -35379 -12933
rect -35424 -12960 -35415 -12942
rect -35388 -12960 -35379 -12942
rect -35361 -12960 -35343 -12933
rect -35316 -12960 -35307 -12933
rect -35874 -12996 -35838 -12987
rect -35874 -13014 -35865 -12996
rect -35847 -13014 -35838 -12996
rect -35820 -13014 -35721 -12987
rect -35703 -13014 -35676 -12987
rect -35658 -13005 -35649 -12987
rect -35631 -13005 -35622 -12987
rect -35658 -13014 -35622 -13005
rect -33426 -12996 -33381 -12987
rect -33426 -13014 -33417 -12996
rect -33390 -13014 -33381 -12996
rect -33363 -13014 -33345 -12987
rect -33318 -13014 -33309 -12987
rect -33876 -13050 -33840 -13041
rect -33876 -13068 -33867 -13050
rect -33849 -13068 -33840 -13050
rect -33822 -13068 -33678 -13041
rect -33660 -13059 -33651 -13041
rect -33633 -13059 -33624 -13041
rect -33660 -13068 -33624 -13059
rect -33426 -13410 -33381 -13401
rect -33426 -13428 -33417 -13410
rect -33390 -13428 -33381 -13410
rect -33363 -13428 -33345 -13401
rect -33318 -13428 -33309 -13401
rect -33876 -13464 -33840 -13455
rect -33876 -13482 -33867 -13464
rect -33849 -13482 -33840 -13464
rect -33822 -13482 -33678 -13455
rect -33660 -13473 -33651 -13455
rect -33633 -13473 -33624 -13455
rect -33660 -13482 -33624 -13473
rect -33426 -13941 -33381 -13932
rect -33426 -13959 -33417 -13941
rect -33390 -13959 -33381 -13941
rect -33363 -13959 -33345 -13932
rect -33318 -13959 -33309 -13932
rect -33876 -13995 -33840 -13986
rect -33876 -14013 -33867 -13995
rect -33849 -14013 -33840 -13995
rect -33822 -14013 -33678 -13986
rect -33660 -14004 -33651 -13986
rect -33633 -14004 -33624 -13986
rect -31455 -13950 -31410 -13941
rect -31455 -13968 -31446 -13950
rect -31419 -13968 -31410 -13950
rect -31392 -13968 -31374 -13941
rect -31347 -13968 -31338 -13941
rect -33660 -14013 -33624 -14004
rect -31905 -14004 -31869 -13995
rect -31905 -14022 -31896 -14004
rect -31878 -14022 -31869 -14004
rect -31851 -14022 -31707 -13995
rect -31689 -14013 -31680 -13995
rect -31662 -14013 -31653 -13995
rect -31689 -14022 -31653 -14013
rect -33426 -14436 -33381 -14427
rect -33426 -14454 -33417 -14436
rect -33390 -14454 -33381 -14436
rect -33363 -14454 -33345 -14427
rect -33318 -14454 -33309 -14427
rect -31455 -14427 -31410 -14418
rect -31455 -14445 -31446 -14427
rect -31419 -14445 -31410 -14427
rect -31392 -14445 -31374 -14418
rect -31347 -14445 -31338 -14418
rect -31905 -14481 -31869 -14472
rect -33876 -14490 -33840 -14481
rect -33876 -14508 -33867 -14490
rect -33849 -14508 -33840 -14490
rect -33822 -14508 -33678 -14481
rect -33660 -14499 -33651 -14481
rect -33633 -14499 -33624 -14481
rect -31905 -14499 -31896 -14481
rect -31878 -14499 -31869 -14481
rect -31851 -14499 -31707 -14472
rect -31689 -14490 -31680 -14472
rect -31662 -14490 -31653 -14472
rect -31689 -14499 -31653 -14490
rect -33660 -14508 -33624 -14499
rect -31455 -14823 -31410 -14814
rect -31455 -14841 -31446 -14823
rect -31419 -14841 -31410 -14823
rect -31392 -14841 -31374 -14814
rect -31347 -14841 -31338 -14814
rect -31905 -14877 -31869 -14868
rect -31905 -14895 -31896 -14877
rect -31878 -14895 -31869 -14877
rect -31851 -14895 -31707 -14868
rect -31689 -14886 -31680 -14868
rect -31662 -14886 -31653 -14868
rect -31689 -14895 -31653 -14886
rect -33426 -14931 -33381 -14922
rect -33426 -14949 -33417 -14931
rect -33390 -14949 -33381 -14931
rect -33363 -14949 -33345 -14922
rect -33318 -14949 -33309 -14922
rect -33876 -14985 -33840 -14976
rect -33876 -15003 -33867 -14985
rect -33849 -15003 -33840 -14985
rect -33822 -15003 -33678 -14976
rect -33660 -14994 -33651 -14976
rect -33633 -14994 -33624 -14976
rect -33660 -15003 -33624 -14994
rect -31455 -15291 -31410 -15282
rect -31455 -15309 -31446 -15291
rect -31419 -15309 -31410 -15291
rect -31392 -15309 -31374 -15282
rect -31347 -15309 -31338 -15282
rect -33426 -15345 -33381 -15336
rect -33426 -15363 -33417 -15345
rect -33390 -15363 -33381 -15345
rect -33363 -15363 -33345 -15336
rect -33318 -15363 -33309 -15336
rect -31905 -15345 -31869 -15336
rect -31905 -15363 -31896 -15345
rect -31878 -15363 -31869 -15345
rect -31851 -15363 -31707 -15336
rect -31689 -15354 -31680 -15336
rect -31662 -15354 -31653 -15336
rect -31689 -15363 -31653 -15354
rect -33876 -15399 -33840 -15390
rect -33876 -15417 -33867 -15399
rect -33849 -15417 -33840 -15399
rect -33822 -15417 -33678 -15390
rect -33660 -15408 -33651 -15390
rect -33633 -15408 -33624 -15390
rect -33660 -15417 -33624 -15408
rect -33426 -15876 -33381 -15867
rect -33426 -15894 -33417 -15876
rect -33390 -15894 -33381 -15876
rect -33363 -15894 -33345 -15867
rect -33318 -15894 -33309 -15867
rect -33876 -15930 -33840 -15921
rect -33876 -15948 -33867 -15930
rect -33849 -15948 -33840 -15930
rect -33822 -15948 -33678 -15921
rect -33660 -15939 -33651 -15921
rect -33633 -15939 -33624 -15921
rect -33660 -15948 -33624 -15939
<< pdiffusion >>
rect -30231 10332 -30168 10341
rect -30231 10296 -30222 10332
rect -30186 10296 -30168 10332
rect -30231 10287 -30168 10296
rect -30231 10260 -30168 10269
rect -30231 10224 -30222 10260
rect -30186 10224 -30168 10260
rect -30231 10215 -30168 10224
rect -30231 10161 -30168 10170
rect -30231 10125 -30222 10161
rect -30186 10125 -30168 10161
rect -30231 10116 -30168 10125
rect -29421 10332 -29358 10341
rect -29421 10296 -29412 10332
rect -29376 10296 -29358 10332
rect -29421 10287 -29358 10296
rect -30231 10089 -30168 10098
rect -30231 10053 -30222 10089
rect -30186 10053 -30168 10089
rect -30231 10044 -30168 10053
rect -30231 9972 -30168 9981
rect -30231 9936 -30222 9972
rect -30186 9936 -30168 9972
rect -30231 9918 -30168 9936
rect -30231 9891 -30168 9900
rect -30231 9855 -30222 9891
rect -30186 9855 -30168 9891
rect -30231 9846 -30168 9855
rect -30231 9810 -30168 9819
rect -30231 9774 -30222 9810
rect -30186 9774 -30168 9810
rect -30231 9756 -30168 9774
rect -30231 9729 -30168 9738
rect -30231 9693 -30222 9729
rect -30186 9693 -30168 9729
rect -30231 9684 -30168 9693
rect -29421 10260 -29358 10269
rect -29421 10224 -29412 10260
rect -29376 10224 -29358 10260
rect -29421 10215 -29358 10224
rect -29421 10161 -29358 10170
rect -29421 10125 -29412 10161
rect -29376 10125 -29358 10161
rect -29421 10116 -29358 10125
rect -28539 10332 -28476 10341
rect -28539 10296 -28530 10332
rect -28494 10296 -28476 10332
rect -28539 10287 -28476 10296
rect -29421 10089 -29358 10098
rect -29421 10053 -29412 10089
rect -29376 10053 -29358 10089
rect -29421 10044 -29358 10053
rect -29421 9972 -29358 9981
rect -29421 9936 -29412 9972
rect -29376 9936 -29358 9972
rect -29421 9918 -29358 9936
rect -29421 9891 -29358 9900
rect -29421 9855 -29412 9891
rect -29376 9855 -29358 9891
rect -29421 9846 -29358 9855
rect -29421 9810 -29358 9819
rect -29421 9774 -29412 9810
rect -29376 9774 -29358 9810
rect -29421 9756 -29358 9774
rect -29421 9729 -29358 9738
rect -29421 9693 -29412 9729
rect -29376 9693 -29358 9729
rect -29421 9684 -29358 9693
rect -28539 10260 -28476 10269
rect -28539 10224 -28530 10260
rect -28494 10224 -28476 10260
rect -28539 10215 -28476 10224
rect -28539 10161 -28476 10170
rect -28539 10125 -28530 10161
rect -28494 10125 -28476 10161
rect -28539 10116 -28476 10125
rect -28539 10089 -28476 10098
rect -28539 10053 -28530 10089
rect -28494 10053 -28476 10089
rect -28539 10044 -28476 10053
rect -28539 9972 -28476 9981
rect -28539 9936 -28530 9972
rect -28494 9936 -28476 9972
rect -28539 9918 -28476 9936
rect -28539 9891 -28476 9900
rect -28539 9855 -28530 9891
rect -28494 9855 -28476 9891
rect -28539 9846 -28476 9855
rect -28539 9810 -28476 9819
rect -28539 9774 -28530 9810
rect -28494 9774 -28476 9810
rect -28539 9756 -28476 9774
rect -28539 9729 -28476 9738
rect -28539 9693 -28530 9729
rect -28494 9693 -28476 9729
rect -28539 9684 -28476 9693
rect -30366 9333 -30330 9342
rect -30366 9315 -30357 9333
rect -30339 9315 -30330 9333
rect -30366 9297 -30330 9315
rect -30312 9324 -30249 9342
rect -30312 9306 -30303 9324
rect -30285 9306 -30249 9324
rect -30312 9297 -30249 9306
rect -30213 9333 -30168 9342
rect -30213 9315 -30204 9333
rect -30186 9315 -30168 9333
rect -30213 9297 -30168 9315
rect -30150 9333 -30114 9342
rect -30150 9315 -30141 9333
rect -30123 9315 -30114 9333
rect -30150 9297 -30114 9315
rect -29916 9351 -29907 9378
rect -29880 9351 -29871 9378
rect -29916 9324 -29871 9351
rect -29853 9369 -29799 9378
rect -29853 9342 -29835 9369
rect -29808 9342 -29799 9369
rect -29853 9324 -29799 9342
rect -29340 9396 -29304 9405
rect -29340 9378 -29331 9396
rect -29313 9378 -29304 9396
rect -29340 9360 -29304 9378
rect -29286 9387 -29223 9405
rect -29286 9369 -29277 9387
rect -29259 9369 -29223 9387
rect -29286 9360 -29223 9369
rect -29187 9396 -29142 9405
rect -29187 9378 -29178 9396
rect -29160 9378 -29142 9396
rect -29187 9360 -29142 9378
rect -29124 9396 -29088 9405
rect -29124 9378 -29115 9396
rect -29097 9378 -29088 9396
rect -29124 9360 -29088 9378
rect -28890 9414 -28881 9441
rect -28854 9414 -28845 9441
rect -28890 9387 -28845 9414
rect -28827 9432 -28773 9441
rect -28827 9405 -28809 9432
rect -28782 9405 -28773 9432
rect -28827 9387 -28773 9405
rect -29700 8973 -29655 8982
rect -29700 8955 -29691 8973
rect -29673 8955 -29655 8973
rect -29700 8937 -29655 8955
rect -29637 8937 -29565 8982
rect -29547 8964 -29520 8982
rect -29547 8946 -29538 8964
rect -29547 8937 -29520 8946
rect -29475 8973 -29439 8982
rect -29475 8955 -29466 8973
rect -29448 8955 -29439 8973
rect -29475 8937 -29439 8955
rect -29421 8964 -29385 8982
rect -29421 8946 -29412 8964
rect -29394 8946 -29385 8964
rect -29421 8937 -29385 8946
rect -30231 8235 -30168 8244
rect -30231 8199 -30222 8235
rect -30186 8199 -30168 8235
rect -30231 8190 -30168 8199
rect -30231 8163 -30168 8172
rect -30231 8127 -30222 8163
rect -30186 8127 -30168 8163
rect -30231 8118 -30168 8127
rect -30231 8064 -30168 8073
rect -30231 8028 -30222 8064
rect -30186 8028 -30168 8064
rect -30231 8019 -30168 8028
rect -29421 8235 -29358 8244
rect -29421 8199 -29412 8235
rect -29376 8199 -29358 8235
rect -29421 8190 -29358 8199
rect -30231 7992 -30168 8001
rect -30231 7956 -30222 7992
rect -30186 7956 -30168 7992
rect -30231 7947 -30168 7956
rect -30231 7875 -30168 7884
rect -30231 7839 -30222 7875
rect -30186 7839 -30168 7875
rect -30231 7821 -30168 7839
rect -30231 7794 -30168 7803
rect -30231 7758 -30222 7794
rect -30186 7758 -30168 7794
rect -30231 7749 -30168 7758
rect -30231 7713 -30168 7722
rect -30231 7677 -30222 7713
rect -30186 7677 -30168 7713
rect -30231 7659 -30168 7677
rect -30231 7632 -30168 7641
rect -30231 7596 -30222 7632
rect -30186 7596 -30168 7632
rect -30231 7587 -30168 7596
rect -29421 8163 -29358 8172
rect -29421 8127 -29412 8163
rect -29376 8127 -29358 8163
rect -29421 8118 -29358 8127
rect -29421 8064 -29358 8073
rect -29421 8028 -29412 8064
rect -29376 8028 -29358 8064
rect -29421 8019 -29358 8028
rect -28539 8235 -28476 8244
rect -28539 8199 -28530 8235
rect -28494 8199 -28476 8235
rect -28539 8190 -28476 8199
rect -29421 7992 -29358 8001
rect -29421 7956 -29412 7992
rect -29376 7956 -29358 7992
rect -29421 7947 -29358 7956
rect -29421 7875 -29358 7884
rect -29421 7839 -29412 7875
rect -29376 7839 -29358 7875
rect -29421 7821 -29358 7839
rect -29421 7794 -29358 7803
rect -29421 7758 -29412 7794
rect -29376 7758 -29358 7794
rect -29421 7749 -29358 7758
rect -29421 7713 -29358 7722
rect -29421 7677 -29412 7713
rect -29376 7677 -29358 7713
rect -29421 7659 -29358 7677
rect -29421 7632 -29358 7641
rect -29421 7596 -29412 7632
rect -29376 7596 -29358 7632
rect -29421 7587 -29358 7596
rect -28539 8163 -28476 8172
rect -28539 8127 -28530 8163
rect -28494 8127 -28476 8163
rect -28539 8118 -28476 8127
rect -28539 8064 -28476 8073
rect -28539 8028 -28530 8064
rect -28494 8028 -28476 8064
rect -28539 8019 -28476 8028
rect -28539 7992 -28476 8001
rect -28539 7956 -28530 7992
rect -28494 7956 -28476 7992
rect -28539 7947 -28476 7956
rect -28539 7875 -28476 7884
rect -28539 7839 -28530 7875
rect -28494 7839 -28476 7875
rect -28539 7821 -28476 7839
rect -28539 7794 -28476 7803
rect -28539 7758 -28530 7794
rect -28494 7758 -28476 7794
rect -28539 7749 -28476 7758
rect -28539 7713 -28476 7722
rect -28539 7677 -28530 7713
rect -28494 7677 -28476 7713
rect -28539 7659 -28476 7677
rect -28539 7632 -28476 7641
rect -28539 7596 -28530 7632
rect -28494 7596 -28476 7632
rect -28539 7587 -28476 7596
rect -30366 7236 -30330 7245
rect -30366 7218 -30357 7236
rect -30339 7218 -30330 7236
rect -30366 7200 -30330 7218
rect -30312 7227 -30249 7245
rect -30312 7209 -30303 7227
rect -30285 7209 -30249 7227
rect -30312 7200 -30249 7209
rect -30213 7236 -30168 7245
rect -30213 7218 -30204 7236
rect -30186 7218 -30168 7236
rect -30213 7200 -30168 7218
rect -30150 7236 -30114 7245
rect -30150 7218 -30141 7236
rect -30123 7218 -30114 7236
rect -30150 7200 -30114 7218
rect -29916 7254 -29907 7281
rect -29880 7254 -29871 7281
rect -29916 7227 -29871 7254
rect -29853 7272 -29799 7281
rect -29853 7245 -29835 7272
rect -29808 7245 -29799 7272
rect -29853 7227 -29799 7245
rect -29340 7299 -29304 7308
rect -29340 7281 -29331 7299
rect -29313 7281 -29304 7299
rect -29340 7263 -29304 7281
rect -29286 7290 -29223 7308
rect -29286 7272 -29277 7290
rect -29259 7272 -29223 7290
rect -29286 7263 -29223 7272
rect -29187 7299 -29142 7308
rect -29187 7281 -29178 7299
rect -29160 7281 -29142 7299
rect -29187 7263 -29142 7281
rect -29124 7299 -29088 7308
rect -29124 7281 -29115 7299
rect -29097 7281 -29088 7299
rect -29124 7263 -29088 7281
rect -28890 7317 -28881 7344
rect -28854 7317 -28845 7344
rect -28890 7290 -28845 7317
rect -28827 7335 -28773 7344
rect -28827 7308 -28809 7335
rect -28782 7308 -28773 7335
rect -28827 7290 -28773 7308
rect -29700 6876 -29655 6885
rect -29700 6858 -29691 6876
rect -29673 6858 -29655 6876
rect -29700 6840 -29655 6858
rect -29637 6840 -29565 6885
rect -29547 6867 -29520 6885
rect -29547 6849 -29538 6867
rect -29547 6840 -29520 6849
rect -29475 6876 -29439 6885
rect -29475 6858 -29466 6876
rect -29448 6858 -29439 6876
rect -29475 6840 -29439 6858
rect -29421 6867 -29385 6885
rect -29421 6849 -29412 6867
rect -29394 6849 -29385 6867
rect -29421 6840 -29385 6849
rect -30231 6120 -30168 6129
rect -30231 6084 -30222 6120
rect -30186 6084 -30168 6120
rect -30231 6075 -30168 6084
rect -30231 6048 -30168 6057
rect -30231 6012 -30222 6048
rect -30186 6012 -30168 6048
rect -30231 6003 -30168 6012
rect -30231 5949 -30168 5958
rect -30231 5913 -30222 5949
rect -30186 5913 -30168 5949
rect -30231 5904 -30168 5913
rect -29421 6120 -29358 6129
rect -29421 6084 -29412 6120
rect -29376 6084 -29358 6120
rect -29421 6075 -29358 6084
rect -30231 5877 -30168 5886
rect -30231 5841 -30222 5877
rect -30186 5841 -30168 5877
rect -30231 5832 -30168 5841
rect -30231 5760 -30168 5769
rect -30231 5724 -30222 5760
rect -30186 5724 -30168 5760
rect -30231 5706 -30168 5724
rect -30231 5679 -30168 5688
rect -30231 5643 -30222 5679
rect -30186 5643 -30168 5679
rect -30231 5634 -30168 5643
rect -30231 5598 -30168 5607
rect -30231 5562 -30222 5598
rect -30186 5562 -30168 5598
rect -30231 5544 -30168 5562
rect -30231 5517 -30168 5526
rect -30231 5481 -30222 5517
rect -30186 5481 -30168 5517
rect -30231 5472 -30168 5481
rect -29421 6048 -29358 6057
rect -29421 6012 -29412 6048
rect -29376 6012 -29358 6048
rect -29421 6003 -29358 6012
rect -29421 5949 -29358 5958
rect -29421 5913 -29412 5949
rect -29376 5913 -29358 5949
rect -29421 5904 -29358 5913
rect -28539 6120 -28476 6129
rect -28539 6084 -28530 6120
rect -28494 6084 -28476 6120
rect -28539 6075 -28476 6084
rect -29421 5877 -29358 5886
rect -29421 5841 -29412 5877
rect -29376 5841 -29358 5877
rect -29421 5832 -29358 5841
rect -29421 5760 -29358 5769
rect -29421 5724 -29412 5760
rect -29376 5724 -29358 5760
rect -29421 5706 -29358 5724
rect -29421 5679 -29358 5688
rect -29421 5643 -29412 5679
rect -29376 5643 -29358 5679
rect -29421 5634 -29358 5643
rect -29421 5598 -29358 5607
rect -29421 5562 -29412 5598
rect -29376 5562 -29358 5598
rect -29421 5544 -29358 5562
rect -29421 5517 -29358 5526
rect -29421 5481 -29412 5517
rect -29376 5481 -29358 5517
rect -29421 5472 -29358 5481
rect -28539 6048 -28476 6057
rect -28539 6012 -28530 6048
rect -28494 6012 -28476 6048
rect -28539 6003 -28476 6012
rect -28539 5949 -28476 5958
rect -28539 5913 -28530 5949
rect -28494 5913 -28476 5949
rect -28539 5904 -28476 5913
rect -28539 5877 -28476 5886
rect -28539 5841 -28530 5877
rect -28494 5841 -28476 5877
rect -28539 5832 -28476 5841
rect -28539 5760 -28476 5769
rect -28539 5724 -28530 5760
rect -28494 5724 -28476 5760
rect -28539 5706 -28476 5724
rect -28539 5679 -28476 5688
rect -28539 5643 -28530 5679
rect -28494 5643 -28476 5679
rect -28539 5634 -28476 5643
rect -28539 5598 -28476 5607
rect -28539 5562 -28530 5598
rect -28494 5562 -28476 5598
rect -28539 5544 -28476 5562
rect -28539 5517 -28476 5526
rect -28539 5481 -28530 5517
rect -28494 5481 -28476 5517
rect -28539 5472 -28476 5481
rect -30366 5121 -30330 5130
rect -30366 5103 -30357 5121
rect -30339 5103 -30330 5121
rect -30366 5085 -30330 5103
rect -30312 5112 -30249 5130
rect -30312 5094 -30303 5112
rect -30285 5094 -30249 5112
rect -30312 5085 -30249 5094
rect -30213 5121 -30168 5130
rect -30213 5103 -30204 5121
rect -30186 5103 -30168 5121
rect -30213 5085 -30168 5103
rect -30150 5121 -30114 5130
rect -30150 5103 -30141 5121
rect -30123 5103 -30114 5121
rect -30150 5085 -30114 5103
rect -29916 5139 -29907 5166
rect -29880 5139 -29871 5166
rect -29916 5112 -29871 5139
rect -29853 5157 -29799 5166
rect -29853 5130 -29835 5157
rect -29808 5130 -29799 5157
rect -29853 5112 -29799 5130
rect -29340 5184 -29304 5193
rect -29340 5166 -29331 5184
rect -29313 5166 -29304 5184
rect -29340 5148 -29304 5166
rect -29286 5175 -29223 5193
rect -29286 5157 -29277 5175
rect -29259 5157 -29223 5175
rect -29286 5148 -29223 5157
rect -29187 5184 -29142 5193
rect -29187 5166 -29178 5184
rect -29160 5166 -29142 5184
rect -29187 5148 -29142 5166
rect -29124 5184 -29088 5193
rect -29124 5166 -29115 5184
rect -29097 5166 -29088 5184
rect -29124 5148 -29088 5166
rect -28890 5202 -28881 5229
rect -28854 5202 -28845 5229
rect -28890 5175 -28845 5202
rect -28827 5220 -28773 5229
rect -28827 5193 -28809 5220
rect -28782 5193 -28773 5220
rect -28827 5175 -28773 5193
rect -29700 4761 -29655 4770
rect -29700 4743 -29691 4761
rect -29673 4743 -29655 4761
rect -29700 4725 -29655 4743
rect -29637 4725 -29565 4770
rect -29547 4752 -29520 4770
rect -29547 4734 -29538 4752
rect -29547 4725 -29520 4734
rect -29475 4761 -29439 4770
rect -29475 4743 -29466 4761
rect -29448 4743 -29439 4761
rect -29475 4725 -29439 4743
rect -29421 4752 -29385 4770
rect -29421 4734 -29412 4752
rect -29394 4734 -29385 4752
rect -29421 4725 -29385 4734
rect -30231 4185 -30168 4194
rect -30231 4149 -30222 4185
rect -30186 4149 -30168 4185
rect -30231 4140 -30168 4149
rect -30231 4113 -30168 4122
rect -30231 4077 -30222 4113
rect -30186 4077 -30168 4113
rect -30231 4068 -30168 4077
rect -30231 4014 -30168 4023
rect -30231 3978 -30222 4014
rect -30186 3978 -30168 4014
rect -30231 3969 -30168 3978
rect -29421 4185 -29358 4194
rect -29421 4149 -29412 4185
rect -29376 4149 -29358 4185
rect -29421 4140 -29358 4149
rect -30231 3942 -30168 3951
rect -30231 3906 -30222 3942
rect -30186 3906 -30168 3942
rect -30231 3897 -30168 3906
rect -30231 3825 -30168 3834
rect -30231 3789 -30222 3825
rect -30186 3789 -30168 3825
rect -30231 3771 -30168 3789
rect -30231 3744 -30168 3753
rect -30231 3708 -30222 3744
rect -30186 3708 -30168 3744
rect -30231 3699 -30168 3708
rect -30231 3663 -30168 3672
rect -30231 3627 -30222 3663
rect -30186 3627 -30168 3663
rect -30231 3609 -30168 3627
rect -30231 3582 -30168 3591
rect -30231 3546 -30222 3582
rect -30186 3546 -30168 3582
rect -30231 3537 -30168 3546
rect -29421 4113 -29358 4122
rect -29421 4077 -29412 4113
rect -29376 4077 -29358 4113
rect -29421 4068 -29358 4077
rect -29421 4014 -29358 4023
rect -29421 3978 -29412 4014
rect -29376 3978 -29358 4014
rect -29421 3969 -29358 3978
rect -28539 4185 -28476 4194
rect -28539 4149 -28530 4185
rect -28494 4149 -28476 4185
rect -28539 4140 -28476 4149
rect -29421 3942 -29358 3951
rect -29421 3906 -29412 3942
rect -29376 3906 -29358 3942
rect -29421 3897 -29358 3906
rect -29421 3825 -29358 3834
rect -29421 3789 -29412 3825
rect -29376 3789 -29358 3825
rect -29421 3771 -29358 3789
rect -29421 3744 -29358 3753
rect -29421 3708 -29412 3744
rect -29376 3708 -29358 3744
rect -29421 3699 -29358 3708
rect -29421 3663 -29358 3672
rect -29421 3627 -29412 3663
rect -29376 3627 -29358 3663
rect -29421 3609 -29358 3627
rect -29421 3582 -29358 3591
rect -29421 3546 -29412 3582
rect -29376 3546 -29358 3582
rect -29421 3537 -29358 3546
rect -28539 4113 -28476 4122
rect -28539 4077 -28530 4113
rect -28494 4077 -28476 4113
rect -28539 4068 -28476 4077
rect -28539 4014 -28476 4023
rect -28539 3978 -28530 4014
rect -28494 3978 -28476 4014
rect -28539 3969 -28476 3978
rect -28539 3942 -28476 3951
rect -28539 3906 -28530 3942
rect -28494 3906 -28476 3942
rect -28539 3897 -28476 3906
rect -28539 3825 -28476 3834
rect -28539 3789 -28530 3825
rect -28494 3789 -28476 3825
rect -28539 3771 -28476 3789
rect -28539 3744 -28476 3753
rect -28539 3708 -28530 3744
rect -28494 3708 -28476 3744
rect -28539 3699 -28476 3708
rect -28539 3663 -28476 3672
rect -28539 3627 -28530 3663
rect -28494 3627 -28476 3663
rect -28539 3609 -28476 3627
rect -28539 3582 -28476 3591
rect -28539 3546 -28530 3582
rect -28494 3546 -28476 3582
rect -28539 3537 -28476 3546
rect -30366 3186 -30330 3195
rect -30366 3168 -30357 3186
rect -30339 3168 -30330 3186
rect -30366 3150 -30330 3168
rect -30312 3177 -30249 3195
rect -30312 3159 -30303 3177
rect -30285 3159 -30249 3177
rect -30312 3150 -30249 3159
rect -30213 3186 -30168 3195
rect -30213 3168 -30204 3186
rect -30186 3168 -30168 3186
rect -30213 3150 -30168 3168
rect -30150 3186 -30114 3195
rect -30150 3168 -30141 3186
rect -30123 3168 -30114 3186
rect -30150 3150 -30114 3168
rect -29916 3204 -29907 3231
rect -29880 3204 -29871 3231
rect -29916 3177 -29871 3204
rect -29853 3222 -29799 3231
rect -29853 3195 -29835 3222
rect -29808 3195 -29799 3222
rect -29853 3177 -29799 3195
rect -29340 3249 -29304 3258
rect -29340 3231 -29331 3249
rect -29313 3231 -29304 3249
rect -29340 3213 -29304 3231
rect -29286 3240 -29223 3258
rect -29286 3222 -29277 3240
rect -29259 3222 -29223 3240
rect -29286 3213 -29223 3222
rect -29187 3249 -29142 3258
rect -29187 3231 -29178 3249
rect -29160 3231 -29142 3249
rect -29187 3213 -29142 3231
rect -29124 3249 -29088 3258
rect -29124 3231 -29115 3249
rect -29097 3231 -29088 3249
rect -29124 3213 -29088 3231
rect -28890 3267 -28881 3294
rect -28854 3267 -28845 3294
rect -28890 3240 -28845 3267
rect -28827 3285 -28773 3294
rect -28827 3258 -28809 3285
rect -28782 3258 -28773 3285
rect -28827 3240 -28773 3258
rect -29700 2826 -29655 2835
rect -29700 2808 -29691 2826
rect -29673 2808 -29655 2826
rect -29700 2790 -29655 2808
rect -29637 2790 -29565 2835
rect -29547 2817 -29520 2835
rect -29547 2799 -29538 2817
rect -29547 2790 -29520 2799
rect -29475 2826 -29439 2835
rect -29475 2808 -29466 2826
rect -29448 2808 -29439 2826
rect -29475 2790 -29439 2808
rect -29421 2817 -29385 2835
rect -29421 2799 -29412 2817
rect -29394 2799 -29385 2817
rect -29421 2790 -29385 2799
rect -29871 495 -29808 504
rect -29871 459 -29862 495
rect -29826 459 -29808 495
rect -29871 450 -29808 459
rect -29871 423 -29808 432
rect -29871 387 -29862 423
rect -29826 387 -29808 423
rect -29871 378 -29808 387
rect -29871 324 -29808 333
rect -29871 288 -29862 324
rect -29826 288 -29808 324
rect -29871 279 -29808 288
rect -29520 369 -29511 396
rect -29484 369 -29475 396
rect -29520 342 -29475 369
rect -29457 387 -29403 396
rect -29457 360 -29439 387
rect -29412 360 -29403 387
rect -29457 342 -29403 360
rect -29871 252 -29808 261
rect -29871 216 -29862 252
rect -29826 216 -29808 252
rect -29871 207 -29808 216
rect -29871 135 -29808 144
rect -29871 99 -29862 135
rect -29826 99 -29808 135
rect -29871 81 -29808 99
rect -29871 54 -29808 63
rect -29871 18 -29862 54
rect -29826 18 -29808 54
rect -29871 9 -29808 18
rect -29871 -27 -29808 -18
rect -29871 -63 -29862 -27
rect -29826 -63 -29808 -27
rect -29871 -81 -29808 -63
rect -29871 -108 -29808 -99
rect -29871 -144 -29862 -108
rect -29826 -144 -29808 -108
rect -29871 -153 -29808 -144
rect -28314 99 -28305 126
rect -28278 99 -28269 126
rect -29151 63 -29142 90
rect -29115 63 -29106 90
rect -29151 36 -29106 63
rect -29088 81 -29034 90
rect -29088 54 -29070 81
rect -29043 54 -29034 81
rect -29088 36 -29034 54
rect -28764 81 -28728 90
rect -28764 63 -28755 81
rect -28737 63 -28728 81
rect -28764 45 -28728 63
rect -28710 72 -28647 90
rect -28710 54 -28701 72
rect -28683 54 -28647 72
rect -28710 45 -28647 54
rect -28611 81 -28566 90
rect -28611 63 -28602 81
rect -28584 63 -28566 81
rect -28611 45 -28566 63
rect -28548 81 -28512 90
rect -28548 63 -28539 81
rect -28521 63 -28512 81
rect -28314 72 -28269 99
rect -28251 117 -28197 126
rect -28251 90 -28233 117
rect -28206 90 -28197 117
rect -28251 72 -28197 90
rect -28548 45 -28512 63
rect -33444 -315 -33435 -288
rect -33408 -315 -33399 -288
rect -33894 -333 -33858 -324
rect -33894 -351 -33885 -333
rect -33867 -351 -33858 -333
rect -33894 -369 -33858 -351
rect -33840 -342 -33777 -324
rect -33840 -360 -33831 -342
rect -33813 -360 -33777 -342
rect -33840 -369 -33777 -360
rect -33741 -333 -33696 -324
rect -33741 -351 -33732 -333
rect -33714 -351 -33696 -333
rect -33741 -369 -33696 -351
rect -33678 -333 -33642 -324
rect -33678 -351 -33669 -333
rect -33651 -351 -33642 -333
rect -33444 -342 -33399 -315
rect -33381 -297 -33327 -288
rect -33381 -324 -33363 -297
rect -33336 -324 -33327 -297
rect -33381 -342 -33327 -324
rect -33678 -369 -33642 -351
rect -29871 -450 -29808 -441
rect -29871 -486 -29862 -450
rect -29826 -486 -29808 -450
rect -29871 -495 -29808 -486
rect -33444 -810 -33435 -783
rect -33408 -810 -33399 -783
rect -33894 -828 -33858 -819
rect -33894 -846 -33885 -828
rect -33867 -846 -33858 -828
rect -33894 -864 -33858 -846
rect -33840 -837 -33777 -819
rect -33840 -855 -33831 -837
rect -33813 -855 -33777 -837
rect -33840 -864 -33777 -855
rect -33741 -828 -33696 -819
rect -33741 -846 -33732 -828
rect -33714 -846 -33696 -828
rect -33741 -864 -33696 -846
rect -33678 -828 -33642 -819
rect -33678 -846 -33669 -828
rect -33651 -846 -33642 -828
rect -33444 -837 -33399 -810
rect -33381 -792 -33327 -783
rect -33381 -819 -33363 -792
rect -33336 -819 -33327 -792
rect -33381 -837 -33327 -819
rect -33678 -864 -33642 -846
rect -34470 -1080 -34425 -1071
rect -34470 -1098 -34461 -1080
rect -34443 -1098 -34425 -1080
rect -34470 -1116 -34425 -1098
rect -34407 -1116 -34335 -1071
rect -34317 -1089 -34290 -1071
rect -34317 -1107 -34308 -1089
rect -34317 -1116 -34290 -1107
rect -34245 -1080 -34209 -1071
rect -34245 -1098 -34236 -1080
rect -34218 -1098 -34209 -1080
rect -34245 -1116 -34209 -1098
rect -34191 -1089 -34155 -1071
rect -34191 -1107 -34182 -1089
rect -34164 -1107 -34155 -1089
rect -34191 -1116 -34155 -1107
rect -33444 -1224 -33435 -1197
rect -33408 -1224 -33399 -1197
rect -33894 -1242 -33858 -1233
rect -33894 -1260 -33885 -1242
rect -33867 -1260 -33858 -1242
rect -33894 -1278 -33858 -1260
rect -33840 -1251 -33777 -1233
rect -33840 -1269 -33831 -1251
rect -33813 -1269 -33777 -1251
rect -33840 -1278 -33777 -1269
rect -33741 -1242 -33696 -1233
rect -33741 -1260 -33732 -1242
rect -33714 -1260 -33696 -1242
rect -33741 -1278 -33696 -1260
rect -33678 -1242 -33642 -1233
rect -33678 -1260 -33669 -1242
rect -33651 -1260 -33642 -1242
rect -33444 -1251 -33399 -1224
rect -33381 -1206 -33327 -1197
rect -33381 -1233 -33363 -1206
rect -33336 -1233 -33327 -1206
rect -33381 -1251 -33327 -1233
rect -33678 -1278 -33642 -1260
rect -33444 -1755 -33435 -1728
rect -33408 -1755 -33399 -1728
rect -33894 -1773 -33858 -1764
rect -33894 -1791 -33885 -1773
rect -33867 -1791 -33858 -1773
rect -33894 -1809 -33858 -1791
rect -33840 -1782 -33777 -1764
rect -33840 -1800 -33831 -1782
rect -33813 -1800 -33777 -1782
rect -33840 -1809 -33777 -1800
rect -33741 -1773 -33696 -1764
rect -33741 -1791 -33732 -1773
rect -33714 -1791 -33696 -1773
rect -33741 -1809 -33696 -1791
rect -33678 -1773 -33642 -1764
rect -33678 -1791 -33669 -1773
rect -33651 -1791 -33642 -1773
rect -33444 -1782 -33399 -1755
rect -33381 -1737 -33327 -1728
rect -33381 -1764 -33363 -1737
rect -33336 -1764 -33327 -1737
rect -33381 -1782 -33327 -1764
rect -33678 -1809 -33642 -1791
rect -33444 -2322 -33435 -2295
rect -33408 -2322 -33399 -2295
rect -33894 -2340 -33858 -2331
rect -33894 -2358 -33885 -2340
rect -33867 -2358 -33858 -2340
rect -33894 -2376 -33858 -2358
rect -33840 -2349 -33777 -2331
rect -33840 -2367 -33831 -2349
rect -33813 -2367 -33777 -2349
rect -33840 -2376 -33777 -2367
rect -33741 -2340 -33696 -2331
rect -33741 -2358 -33732 -2340
rect -33714 -2358 -33696 -2340
rect -33741 -2376 -33696 -2358
rect -33678 -2340 -33642 -2331
rect -33678 -2358 -33669 -2340
rect -33651 -2358 -33642 -2340
rect -33444 -2349 -33399 -2322
rect -33381 -2304 -33327 -2295
rect -33381 -2331 -33363 -2304
rect -33336 -2331 -33327 -2304
rect -33381 -2349 -33327 -2331
rect -33678 -2376 -33642 -2358
rect -33444 -2817 -33435 -2790
rect -33408 -2817 -33399 -2790
rect -33894 -2835 -33858 -2826
rect -33894 -2853 -33885 -2835
rect -33867 -2853 -33858 -2835
rect -33894 -2871 -33858 -2853
rect -33840 -2844 -33777 -2826
rect -33840 -2862 -33831 -2844
rect -33813 -2862 -33777 -2844
rect -33840 -2871 -33777 -2862
rect -33741 -2835 -33696 -2826
rect -33741 -2853 -33732 -2835
rect -33714 -2853 -33696 -2835
rect -33741 -2871 -33696 -2853
rect -33678 -2835 -33642 -2826
rect -33678 -2853 -33669 -2835
rect -33651 -2853 -33642 -2835
rect -33444 -2844 -33399 -2817
rect -33381 -2799 -33327 -2790
rect -33381 -2826 -33363 -2799
rect -33336 -2826 -33327 -2799
rect -33381 -2844 -33327 -2826
rect -33678 -2871 -33642 -2853
rect -33444 -3231 -33435 -3204
rect -33408 -3231 -33399 -3204
rect -33894 -3249 -33858 -3240
rect -33894 -3267 -33885 -3249
rect -33867 -3267 -33858 -3249
rect -33894 -3285 -33858 -3267
rect -33840 -3258 -33777 -3240
rect -33840 -3276 -33831 -3258
rect -33813 -3276 -33777 -3258
rect -33840 -3285 -33777 -3276
rect -33741 -3249 -33696 -3240
rect -33741 -3267 -33732 -3249
rect -33714 -3267 -33696 -3249
rect -33741 -3285 -33696 -3267
rect -33678 -3249 -33642 -3240
rect -33678 -3267 -33669 -3249
rect -33651 -3267 -33642 -3249
rect -33444 -3258 -33399 -3231
rect -33381 -3213 -33327 -3204
rect -33381 -3240 -33363 -3213
rect -33336 -3240 -33327 -3213
rect -33381 -3258 -33327 -3240
rect -33678 -3285 -33642 -3267
rect -33444 -3762 -33435 -3735
rect -33408 -3762 -33399 -3735
rect -33894 -3780 -33858 -3771
rect -33894 -3798 -33885 -3780
rect -33867 -3798 -33858 -3780
rect -33894 -3816 -33858 -3798
rect -33840 -3789 -33777 -3771
rect -33840 -3807 -33831 -3789
rect -33813 -3807 -33777 -3789
rect -33840 -3816 -33777 -3807
rect -33741 -3780 -33696 -3771
rect -33741 -3798 -33732 -3780
rect -33714 -3798 -33696 -3780
rect -33741 -3816 -33696 -3798
rect -33678 -3780 -33642 -3771
rect -33678 -3798 -33669 -3780
rect -33651 -3798 -33642 -3780
rect -33444 -3789 -33399 -3762
rect -33381 -3744 -33327 -3735
rect -33381 -3771 -33363 -3744
rect -33336 -3771 -33327 -3744
rect -33381 -3789 -33327 -3771
rect -33678 -3816 -33642 -3798
rect -33426 -8172 -33417 -8145
rect -33390 -8172 -33381 -8145
rect -33876 -8190 -33840 -8181
rect -33876 -8208 -33867 -8190
rect -33849 -8208 -33840 -8190
rect -33876 -8226 -33840 -8208
rect -33822 -8199 -33759 -8181
rect -33822 -8217 -33813 -8199
rect -33795 -8217 -33759 -8199
rect -33822 -8226 -33759 -8217
rect -33723 -8190 -33678 -8181
rect -33723 -8208 -33714 -8190
rect -33696 -8208 -33678 -8190
rect -33723 -8226 -33678 -8208
rect -33660 -8190 -33624 -8181
rect -33660 -8208 -33651 -8190
rect -33633 -8208 -33624 -8190
rect -33426 -8199 -33381 -8172
rect -33363 -8154 -33309 -8145
rect -33363 -8181 -33345 -8154
rect -33318 -8181 -33309 -8154
rect -33363 -8199 -33309 -8181
rect -33660 -8226 -33624 -8208
rect -29871 -522 -29808 -513
rect -29871 -558 -29862 -522
rect -29826 -558 -29808 -522
rect -29871 -567 -29808 -558
rect -29871 -621 -29808 -612
rect -29871 -657 -29862 -621
rect -29826 -657 -29808 -621
rect -29871 -666 -29808 -657
rect -29520 -576 -29511 -549
rect -29484 -576 -29475 -549
rect -29520 -603 -29475 -576
rect -29457 -558 -29403 -549
rect -29457 -585 -29439 -558
rect -29412 -585 -29403 -558
rect -29457 -603 -29403 -585
rect -29871 -693 -29808 -684
rect -29871 -729 -29862 -693
rect -29826 -729 -29808 -693
rect -28386 -711 -28377 -684
rect -28350 -711 -28341 -684
rect -29871 -738 -29808 -729
rect -29871 -810 -29808 -801
rect -29871 -846 -29862 -810
rect -29826 -846 -29808 -810
rect -29871 -864 -29808 -846
rect -29871 -891 -29808 -882
rect -29871 -927 -29862 -891
rect -29826 -927 -29808 -891
rect -29169 -747 -29160 -720
rect -29133 -747 -29124 -720
rect -29169 -774 -29124 -747
rect -29106 -729 -29052 -720
rect -29106 -756 -29088 -729
rect -29061 -756 -29052 -729
rect -29106 -774 -29052 -756
rect -28836 -729 -28800 -720
rect -28836 -747 -28827 -729
rect -28809 -747 -28800 -729
rect -28836 -765 -28800 -747
rect -28782 -738 -28719 -720
rect -28782 -756 -28773 -738
rect -28755 -756 -28719 -738
rect -28782 -765 -28719 -756
rect -28683 -729 -28638 -720
rect -28683 -747 -28674 -729
rect -28656 -747 -28638 -729
rect -28683 -765 -28638 -747
rect -28620 -729 -28584 -720
rect -28620 -747 -28611 -729
rect -28593 -747 -28584 -729
rect -28386 -738 -28341 -711
rect -28323 -693 -28269 -684
rect -28323 -720 -28305 -693
rect -28278 -720 -28269 -693
rect -28323 -738 -28269 -720
rect -28008 -729 -27972 -720
rect -28620 -765 -28584 -747
rect -28008 -747 -27999 -729
rect -27981 -747 -27972 -729
rect -28008 -765 -27972 -747
rect -27954 -738 -27891 -720
rect -27954 -756 -27945 -738
rect -27927 -756 -27891 -738
rect -27954 -765 -27891 -756
rect -27558 -711 -27549 -684
rect -27522 -711 -27513 -684
rect -27855 -729 -27810 -720
rect -27855 -747 -27846 -729
rect -27828 -747 -27810 -729
rect -27855 -765 -27810 -747
rect -27792 -729 -27756 -720
rect -27792 -747 -27783 -729
rect -27765 -747 -27756 -729
rect -27558 -738 -27513 -711
rect -27495 -693 -27441 -684
rect -27495 -720 -27477 -693
rect -27450 -720 -27441 -693
rect -27495 -738 -27441 -720
rect -27135 -738 -27090 -729
rect -27792 -765 -27756 -747
rect -27135 -756 -27126 -738
rect -27108 -756 -27090 -738
rect -27135 -774 -27090 -756
rect -27072 -774 -27036 -729
rect -27018 -774 -27000 -729
rect -26982 -774 -26910 -729
rect -26892 -774 -26820 -729
rect -26802 -747 -26775 -729
rect -26802 -765 -26793 -747
rect -26802 -774 -26775 -765
rect -26730 -738 -26694 -729
rect -26730 -756 -26721 -738
rect -26703 -756 -26694 -738
rect -26730 -774 -26694 -756
rect -26676 -747 -26640 -729
rect -26676 -765 -26667 -747
rect -26649 -765 -26640 -747
rect -26676 -774 -26640 -765
rect -29871 -936 -29808 -927
rect -29871 -972 -29808 -963
rect -29871 -1008 -29862 -972
rect -29826 -1008 -29808 -972
rect -29871 -1026 -29808 -1008
rect -29871 -1053 -29808 -1044
rect -29871 -1089 -29862 -1053
rect -29826 -1089 -29808 -1053
rect -29871 -1098 -29808 -1089
rect -29871 -1467 -29808 -1458
rect -29871 -1503 -29862 -1467
rect -29826 -1503 -29808 -1467
rect -29871 -1512 -29808 -1503
rect -29871 -1539 -29808 -1530
rect -29871 -1575 -29862 -1539
rect -29826 -1575 -29808 -1539
rect -29871 -1584 -29808 -1575
rect -29871 -1638 -29808 -1629
rect -29871 -1674 -29862 -1638
rect -29826 -1674 -29808 -1638
rect -29871 -1683 -29808 -1674
rect -28683 -1503 -28638 -1494
rect -28683 -1530 -28674 -1503
rect -28647 -1530 -28638 -1503
rect -28683 -1548 -28638 -1530
rect -28620 -1512 -28575 -1494
rect -28620 -1539 -28611 -1512
rect -28584 -1539 -28575 -1512
rect -28620 -1548 -28575 -1539
rect -28557 -1503 -28512 -1494
rect -28557 -1530 -28548 -1503
rect -28521 -1530 -28512 -1503
rect -28557 -1548 -28512 -1530
rect -28494 -1512 -28440 -1494
rect -28494 -1539 -28485 -1512
rect -28458 -1539 -28440 -1512
rect -28494 -1548 -28440 -1539
rect -28422 -1503 -28368 -1494
rect -28422 -1530 -28404 -1503
rect -28377 -1530 -28368 -1503
rect -28422 -1548 -28368 -1530
rect -28350 -1512 -28305 -1494
rect -28350 -1539 -28341 -1512
rect -28314 -1539 -28305 -1512
rect -28350 -1548 -28305 -1539
rect -28287 -1503 -28242 -1494
rect -28287 -1530 -28278 -1503
rect -28251 -1530 -28242 -1503
rect -28287 -1548 -28242 -1530
rect -28224 -1512 -28179 -1494
rect -28224 -1539 -28215 -1512
rect -28188 -1539 -28179 -1512
rect -28224 -1548 -28179 -1539
rect -28161 -1503 -28107 -1494
rect -28161 -1530 -28152 -1503
rect -28125 -1530 -28107 -1503
rect -28161 -1548 -28107 -1530
rect -28089 -1512 -27954 -1494
rect -28089 -1539 -28080 -1512
rect -28053 -1539 -27954 -1512
rect -28089 -1548 -27954 -1539
rect -27900 -1521 -27882 -1494
rect -27855 -1521 -27846 -1494
rect -27900 -1548 -27846 -1521
rect -27828 -1512 -27783 -1494
rect -27828 -1539 -27819 -1512
rect -27792 -1539 -27783 -1512
rect -27828 -1548 -27783 -1539
rect -29520 -1593 -29511 -1566
rect -29484 -1593 -29475 -1566
rect -29520 -1620 -29475 -1593
rect -29457 -1575 -29403 -1566
rect -29457 -1602 -29439 -1575
rect -29412 -1602 -29403 -1575
rect -29457 -1620 -29403 -1602
rect -29187 -1593 -29178 -1566
rect -29151 -1593 -29142 -1566
rect -29187 -1620 -29142 -1593
rect -29124 -1575 -29070 -1566
rect -29124 -1602 -29106 -1575
rect -29079 -1602 -29070 -1575
rect -29124 -1620 -29070 -1602
rect -29871 -1710 -29808 -1701
rect -29871 -1746 -29862 -1710
rect -29826 -1746 -29808 -1710
rect -29871 -1755 -29808 -1746
rect -29871 -1827 -29808 -1818
rect -29871 -1863 -29862 -1827
rect -29826 -1863 -29808 -1827
rect -29871 -1881 -29808 -1863
rect -29871 -1908 -29808 -1899
rect -29871 -1944 -29862 -1908
rect -29826 -1944 -29808 -1908
rect -29871 -1953 -29808 -1944
rect -29871 -1989 -29808 -1980
rect -29871 -2025 -29862 -1989
rect -29826 -2025 -29808 -1989
rect -29871 -2043 -29808 -2025
rect -29871 -2070 -29808 -2061
rect -29871 -2106 -29862 -2070
rect -29826 -2106 -29808 -2070
rect -29871 -2115 -29808 -2106
rect -29871 -2763 -29808 -2754
rect -29871 -2799 -29862 -2763
rect -29826 -2799 -29808 -2763
rect -29871 -2808 -29808 -2799
rect -29871 -2835 -29808 -2826
rect -29871 -2871 -29862 -2835
rect -29826 -2871 -29808 -2835
rect -29871 -2880 -29808 -2871
rect -29871 -2934 -29808 -2925
rect -29871 -2970 -29862 -2934
rect -29826 -2970 -29808 -2934
rect -29871 -2979 -29808 -2970
rect -28836 -2799 -28791 -2790
rect -28836 -2826 -28827 -2799
rect -28800 -2826 -28791 -2799
rect -28836 -2844 -28791 -2826
rect -28773 -2808 -28728 -2790
rect -28773 -2835 -28764 -2808
rect -28737 -2835 -28728 -2808
rect -28773 -2844 -28728 -2835
rect -28710 -2799 -28665 -2790
rect -28710 -2826 -28701 -2799
rect -28674 -2826 -28665 -2799
rect -28710 -2844 -28665 -2826
rect -28647 -2808 -28593 -2790
rect -28647 -2835 -28638 -2808
rect -28611 -2835 -28593 -2808
rect -28647 -2844 -28593 -2835
rect -28575 -2799 -28521 -2790
rect -28575 -2826 -28557 -2799
rect -28530 -2826 -28521 -2799
rect -28575 -2844 -28521 -2826
rect -28503 -2808 -28458 -2790
rect -28503 -2835 -28494 -2808
rect -28467 -2835 -28458 -2808
rect -28503 -2844 -28458 -2835
rect -28440 -2799 -28395 -2790
rect -28440 -2826 -28431 -2799
rect -28404 -2826 -28395 -2799
rect -28440 -2844 -28395 -2826
rect -28377 -2808 -28332 -2790
rect -28377 -2835 -28368 -2808
rect -28341 -2835 -28332 -2808
rect -28377 -2844 -28332 -2835
rect -28314 -2799 -28260 -2790
rect -28314 -2826 -28305 -2799
rect -28278 -2826 -28260 -2799
rect -28314 -2844 -28260 -2826
rect -28242 -2808 -28107 -2790
rect -28242 -2835 -28233 -2808
rect -28206 -2835 -28107 -2808
rect -28242 -2844 -28107 -2835
rect -28053 -2817 -28035 -2790
rect -28008 -2817 -27999 -2790
rect -28053 -2844 -27999 -2817
rect -27981 -2808 -27936 -2790
rect -27981 -2835 -27972 -2808
rect -27945 -2835 -27936 -2808
rect -27981 -2844 -27936 -2835
rect -29520 -2889 -29511 -2862
rect -29484 -2889 -29475 -2862
rect -29520 -2916 -29475 -2889
rect -29457 -2871 -29403 -2862
rect -29457 -2898 -29439 -2871
rect -29412 -2898 -29403 -2871
rect -29457 -2916 -29403 -2898
rect -29241 -2889 -29232 -2862
rect -29205 -2889 -29196 -2862
rect -29241 -2916 -29196 -2889
rect -29178 -2871 -29124 -2862
rect -29178 -2898 -29160 -2871
rect -29133 -2898 -29124 -2871
rect -29178 -2916 -29124 -2898
rect -29871 -3006 -29808 -2997
rect -29871 -3042 -29862 -3006
rect -29826 -3042 -29808 -3006
rect -29871 -3051 -29808 -3042
rect -29871 -3123 -29808 -3114
rect -29871 -3159 -29862 -3123
rect -29826 -3159 -29808 -3123
rect -29871 -3177 -29808 -3159
rect -29871 -3204 -29808 -3195
rect -29871 -3240 -29862 -3204
rect -29826 -3240 -29808 -3204
rect -29871 -3249 -29808 -3240
rect -29871 -3285 -29808 -3276
rect -29871 -3321 -29862 -3285
rect -29826 -3321 -29808 -3285
rect -29871 -3339 -29808 -3321
rect -29871 -3366 -29808 -3357
rect -29871 -3402 -29862 -3366
rect -29826 -3402 -29808 -3366
rect -29871 -3411 -29808 -3402
rect -29871 -3834 -29808 -3825
rect -29871 -3870 -29862 -3834
rect -29826 -3870 -29808 -3834
rect -29871 -3879 -29808 -3870
rect -29871 -3906 -29808 -3897
rect -29871 -3942 -29862 -3906
rect -29826 -3942 -29808 -3906
rect -29871 -3951 -29808 -3942
rect -29871 -4005 -29808 -3996
rect -29871 -4041 -29862 -4005
rect -29826 -4041 -29808 -4005
rect -29871 -4050 -29808 -4041
rect -29520 -3960 -29511 -3933
rect -29484 -3960 -29475 -3933
rect -29520 -3987 -29475 -3960
rect -29457 -3942 -29403 -3933
rect -29457 -3969 -29439 -3942
rect -29412 -3969 -29403 -3942
rect -29457 -3987 -29403 -3969
rect -29871 -4077 -29808 -4068
rect -29871 -4113 -29862 -4077
rect -29826 -4113 -29808 -4077
rect -29871 -4122 -29808 -4113
rect -29871 -4194 -29808 -4185
rect -29871 -4230 -29862 -4194
rect -29826 -4230 -29808 -4194
rect -29871 -4248 -29808 -4230
rect -29871 -4275 -29808 -4266
rect -29871 -4311 -29862 -4275
rect -29826 -4311 -29808 -4275
rect -29871 -4320 -29808 -4311
rect -29871 -4356 -29808 -4347
rect -29871 -4392 -29862 -4356
rect -29826 -4392 -29808 -4356
rect -29871 -4410 -29808 -4392
rect -29871 -4437 -29808 -4428
rect -29871 -4473 -29862 -4437
rect -29826 -4473 -29808 -4437
rect -29871 -4482 -29808 -4473
rect -28314 -4230 -28305 -4203
rect -28278 -4230 -28269 -4203
rect -29151 -4266 -29142 -4239
rect -29115 -4266 -29106 -4239
rect -29151 -4293 -29106 -4266
rect -29088 -4248 -29034 -4239
rect -29088 -4275 -29070 -4248
rect -29043 -4275 -29034 -4248
rect -29088 -4293 -29034 -4275
rect -28764 -4248 -28728 -4239
rect -28764 -4266 -28755 -4248
rect -28737 -4266 -28728 -4248
rect -28764 -4284 -28728 -4266
rect -28710 -4257 -28647 -4239
rect -28710 -4275 -28701 -4257
rect -28683 -4275 -28647 -4257
rect -28710 -4284 -28647 -4275
rect -28611 -4248 -28566 -4239
rect -28611 -4266 -28602 -4248
rect -28584 -4266 -28566 -4248
rect -28611 -4284 -28566 -4266
rect -28548 -4248 -28512 -4239
rect -28548 -4266 -28539 -4248
rect -28521 -4266 -28512 -4248
rect -28314 -4257 -28269 -4230
rect -28251 -4212 -28197 -4203
rect -28251 -4239 -28233 -4212
rect -28206 -4239 -28197 -4212
rect -28251 -4257 -28197 -4239
rect -28548 -4284 -28512 -4266
rect -29871 -4779 -29808 -4770
rect -29871 -4815 -29862 -4779
rect -29826 -4815 -29808 -4779
rect -29871 -4824 -29808 -4815
rect -29871 -4851 -29808 -4842
rect -29871 -4887 -29862 -4851
rect -29826 -4887 -29808 -4851
rect -29871 -4896 -29808 -4887
rect -29871 -4950 -29808 -4941
rect -29871 -4986 -29862 -4950
rect -29826 -4986 -29808 -4950
rect -29871 -4995 -29808 -4986
rect -29520 -4905 -29511 -4878
rect -29484 -4905 -29475 -4878
rect -29520 -4932 -29475 -4905
rect -29457 -4887 -29403 -4878
rect -29457 -4914 -29439 -4887
rect -29412 -4914 -29403 -4887
rect -29457 -4932 -29403 -4914
rect -29871 -5022 -29808 -5013
rect -29871 -5058 -29862 -5022
rect -29826 -5058 -29808 -5022
rect -28386 -5040 -28377 -5013
rect -28350 -5040 -28341 -5013
rect -29871 -5067 -29808 -5058
rect -29871 -5139 -29808 -5130
rect -29871 -5175 -29862 -5139
rect -29826 -5175 -29808 -5139
rect -29871 -5193 -29808 -5175
rect -29871 -5220 -29808 -5211
rect -29871 -5256 -29862 -5220
rect -29826 -5256 -29808 -5220
rect -29169 -5076 -29160 -5049
rect -29133 -5076 -29124 -5049
rect -29169 -5103 -29124 -5076
rect -29106 -5058 -29052 -5049
rect -29106 -5085 -29088 -5058
rect -29061 -5085 -29052 -5058
rect -29106 -5103 -29052 -5085
rect -28836 -5058 -28800 -5049
rect -28836 -5076 -28827 -5058
rect -28809 -5076 -28800 -5058
rect -28836 -5094 -28800 -5076
rect -28782 -5067 -28719 -5049
rect -28782 -5085 -28773 -5067
rect -28755 -5085 -28719 -5067
rect -28782 -5094 -28719 -5085
rect -28683 -5058 -28638 -5049
rect -28683 -5076 -28674 -5058
rect -28656 -5076 -28638 -5058
rect -28683 -5094 -28638 -5076
rect -28620 -5058 -28584 -5049
rect -28620 -5076 -28611 -5058
rect -28593 -5076 -28584 -5058
rect -28386 -5067 -28341 -5040
rect -28323 -5022 -28269 -5013
rect -28323 -5049 -28305 -5022
rect -28278 -5049 -28269 -5022
rect -28323 -5067 -28269 -5049
rect -28008 -5058 -27972 -5049
rect -28620 -5094 -28584 -5076
rect -28008 -5076 -27999 -5058
rect -27981 -5076 -27972 -5058
rect -28008 -5094 -27972 -5076
rect -27954 -5067 -27891 -5049
rect -27954 -5085 -27945 -5067
rect -27927 -5085 -27891 -5067
rect -27954 -5094 -27891 -5085
rect -27558 -5040 -27549 -5013
rect -27522 -5040 -27513 -5013
rect -27855 -5058 -27810 -5049
rect -27855 -5076 -27846 -5058
rect -27828 -5076 -27810 -5058
rect -27855 -5094 -27810 -5076
rect -27792 -5058 -27756 -5049
rect -27792 -5076 -27783 -5058
rect -27765 -5076 -27756 -5058
rect -27558 -5067 -27513 -5040
rect -27495 -5022 -27441 -5013
rect -27495 -5049 -27477 -5022
rect -27450 -5049 -27441 -5022
rect -27495 -5067 -27441 -5049
rect -27135 -5067 -27090 -5058
rect -27792 -5094 -27756 -5076
rect -27135 -5085 -27126 -5067
rect -27108 -5085 -27090 -5067
rect -27135 -5103 -27090 -5085
rect -27072 -5103 -27036 -5058
rect -27018 -5103 -27000 -5058
rect -26982 -5103 -26910 -5058
rect -26892 -5103 -26820 -5058
rect -26802 -5076 -26775 -5058
rect -26802 -5094 -26793 -5076
rect -26802 -5103 -26775 -5094
rect -26730 -5067 -26694 -5058
rect -26730 -5085 -26721 -5067
rect -26703 -5085 -26694 -5067
rect -26730 -5103 -26694 -5085
rect -26676 -5076 -26640 -5058
rect -26676 -5094 -26667 -5076
rect -26649 -5094 -26640 -5076
rect -26676 -5103 -26640 -5094
rect -29871 -5265 -29808 -5256
rect -29871 -5301 -29808 -5292
rect -29871 -5337 -29862 -5301
rect -29826 -5337 -29808 -5301
rect -29871 -5355 -29808 -5337
rect -29871 -5382 -29808 -5373
rect -29871 -5418 -29862 -5382
rect -29826 -5418 -29808 -5382
rect -29871 -5427 -29808 -5418
rect -29871 -5796 -29808 -5787
rect -29871 -5832 -29862 -5796
rect -29826 -5832 -29808 -5796
rect -29871 -5841 -29808 -5832
rect -29871 -5868 -29808 -5859
rect -29871 -5904 -29862 -5868
rect -29826 -5904 -29808 -5868
rect -29871 -5913 -29808 -5904
rect -29871 -5967 -29808 -5958
rect -29871 -6003 -29862 -5967
rect -29826 -6003 -29808 -5967
rect -29871 -6012 -29808 -6003
rect -28683 -5832 -28638 -5823
rect -28683 -5859 -28674 -5832
rect -28647 -5859 -28638 -5832
rect -28683 -5877 -28638 -5859
rect -28620 -5841 -28575 -5823
rect -28620 -5868 -28611 -5841
rect -28584 -5868 -28575 -5841
rect -28620 -5877 -28575 -5868
rect -28557 -5832 -28512 -5823
rect -28557 -5859 -28548 -5832
rect -28521 -5859 -28512 -5832
rect -28557 -5877 -28512 -5859
rect -28494 -5841 -28440 -5823
rect -28494 -5868 -28485 -5841
rect -28458 -5868 -28440 -5841
rect -28494 -5877 -28440 -5868
rect -28422 -5832 -28368 -5823
rect -28422 -5859 -28404 -5832
rect -28377 -5859 -28368 -5832
rect -28422 -5877 -28368 -5859
rect -28350 -5841 -28305 -5823
rect -28350 -5868 -28341 -5841
rect -28314 -5868 -28305 -5841
rect -28350 -5877 -28305 -5868
rect -28287 -5832 -28242 -5823
rect -28287 -5859 -28278 -5832
rect -28251 -5859 -28242 -5832
rect -28287 -5877 -28242 -5859
rect -28224 -5841 -28179 -5823
rect -28224 -5868 -28215 -5841
rect -28188 -5868 -28179 -5841
rect -28224 -5877 -28179 -5868
rect -28161 -5832 -28107 -5823
rect -28161 -5859 -28152 -5832
rect -28125 -5859 -28107 -5832
rect -28161 -5877 -28107 -5859
rect -28089 -5841 -27954 -5823
rect -28089 -5868 -28080 -5841
rect -28053 -5868 -27954 -5841
rect -28089 -5877 -27954 -5868
rect -27900 -5850 -27882 -5823
rect -27855 -5850 -27846 -5823
rect -27900 -5877 -27846 -5850
rect -27828 -5841 -27783 -5823
rect -27828 -5868 -27819 -5841
rect -27792 -5868 -27783 -5841
rect -27828 -5877 -27783 -5868
rect -29520 -5922 -29511 -5895
rect -29484 -5922 -29475 -5895
rect -29520 -5949 -29475 -5922
rect -29457 -5904 -29403 -5895
rect -29457 -5931 -29439 -5904
rect -29412 -5931 -29403 -5904
rect -29457 -5949 -29403 -5931
rect -29187 -5922 -29178 -5895
rect -29151 -5922 -29142 -5895
rect -29187 -5949 -29142 -5922
rect -29124 -5904 -29070 -5895
rect -29124 -5931 -29106 -5904
rect -29079 -5931 -29070 -5904
rect -29124 -5949 -29070 -5931
rect -29871 -6039 -29808 -6030
rect -29871 -6075 -29862 -6039
rect -29826 -6075 -29808 -6039
rect -29871 -6084 -29808 -6075
rect -29871 -6156 -29808 -6147
rect -29871 -6192 -29862 -6156
rect -29826 -6192 -29808 -6156
rect -29871 -6210 -29808 -6192
rect -29871 -6237 -29808 -6228
rect -29871 -6273 -29862 -6237
rect -29826 -6273 -29808 -6237
rect -29871 -6282 -29808 -6273
rect -29871 -6318 -29808 -6309
rect -29871 -6354 -29862 -6318
rect -29826 -6354 -29808 -6318
rect -29871 -6372 -29808 -6354
rect -29871 -6399 -29808 -6390
rect -29871 -6435 -29862 -6399
rect -29826 -6435 -29808 -6399
rect -29871 -6444 -29808 -6435
rect -33426 -8667 -33417 -8640
rect -33390 -8667 -33381 -8640
rect -33876 -8685 -33840 -8676
rect -33876 -8703 -33867 -8685
rect -33849 -8703 -33840 -8685
rect -33876 -8721 -33840 -8703
rect -33822 -8694 -33759 -8676
rect -33822 -8712 -33813 -8694
rect -33795 -8712 -33759 -8694
rect -33822 -8721 -33759 -8712
rect -33723 -8685 -33678 -8676
rect -33723 -8703 -33714 -8685
rect -33696 -8703 -33678 -8685
rect -33723 -8721 -33678 -8703
rect -33660 -8685 -33624 -8676
rect -33660 -8703 -33651 -8685
rect -33633 -8703 -33624 -8685
rect -33426 -8694 -33381 -8667
rect -33363 -8649 -33309 -8640
rect -33363 -8676 -33345 -8649
rect -33318 -8676 -33309 -8649
rect -33363 -8694 -33309 -8676
rect -33660 -8721 -33624 -8703
rect -33426 -9081 -33417 -9054
rect -33390 -9081 -33381 -9054
rect -33876 -9099 -33840 -9090
rect -33876 -9117 -33867 -9099
rect -33849 -9117 -33840 -9099
rect -33876 -9135 -33840 -9117
rect -33822 -9108 -33759 -9090
rect -33822 -9126 -33813 -9108
rect -33795 -9126 -33759 -9108
rect -33822 -9135 -33759 -9126
rect -33723 -9099 -33678 -9090
rect -33723 -9117 -33714 -9099
rect -33696 -9117 -33678 -9099
rect -33723 -9135 -33678 -9117
rect -33660 -9099 -33624 -9090
rect -33660 -9117 -33651 -9099
rect -33633 -9117 -33624 -9099
rect -33426 -9108 -33381 -9081
rect -33363 -9063 -33309 -9054
rect -33363 -9090 -33345 -9063
rect -33318 -9090 -33309 -9063
rect -33363 -9108 -33309 -9090
rect -33660 -9135 -33624 -9117
rect -33426 -9612 -33417 -9585
rect -33390 -9612 -33381 -9585
rect -33876 -9630 -33840 -9621
rect -33876 -9648 -33867 -9630
rect -33849 -9648 -33840 -9630
rect -33876 -9666 -33840 -9648
rect -33822 -9639 -33759 -9621
rect -33822 -9657 -33813 -9639
rect -33795 -9657 -33759 -9639
rect -33822 -9666 -33759 -9657
rect -33723 -9630 -33678 -9621
rect -33723 -9648 -33714 -9630
rect -33696 -9648 -33678 -9630
rect -33723 -9666 -33678 -9648
rect -33660 -9630 -33624 -9621
rect -33660 -9648 -33651 -9630
rect -33633 -9648 -33624 -9630
rect -33426 -9639 -33381 -9612
rect -33363 -9594 -33309 -9585
rect -33363 -9621 -33345 -9594
rect -33318 -9621 -33309 -9594
rect -33363 -9639 -33309 -9621
rect -33660 -9666 -33624 -9648
rect -33426 -10089 -33417 -10062
rect -33390 -10089 -33381 -10062
rect -33876 -10107 -33840 -10098
rect -33876 -10125 -33867 -10107
rect -33849 -10125 -33840 -10107
rect -33876 -10143 -33840 -10125
rect -33822 -10116 -33759 -10098
rect -33822 -10134 -33813 -10116
rect -33795 -10134 -33759 -10116
rect -33822 -10143 -33759 -10134
rect -33723 -10107 -33678 -10098
rect -33723 -10125 -33714 -10107
rect -33696 -10125 -33678 -10107
rect -33723 -10143 -33678 -10125
rect -33660 -10107 -33624 -10098
rect -33660 -10125 -33651 -10107
rect -33633 -10125 -33624 -10107
rect -33426 -10116 -33381 -10089
rect -33363 -10071 -33309 -10062
rect -33363 -10098 -33345 -10071
rect -33318 -10098 -33309 -10071
rect -33363 -10116 -33309 -10098
rect -33660 -10143 -33624 -10125
rect -33426 -10584 -33417 -10557
rect -33390 -10584 -33381 -10557
rect -33876 -10602 -33840 -10593
rect -33876 -10620 -33867 -10602
rect -33849 -10620 -33840 -10602
rect -33876 -10638 -33840 -10620
rect -33822 -10611 -33759 -10593
rect -33822 -10629 -33813 -10611
rect -33795 -10629 -33759 -10611
rect -33822 -10638 -33759 -10629
rect -33723 -10602 -33678 -10593
rect -33723 -10620 -33714 -10602
rect -33696 -10620 -33678 -10602
rect -33723 -10638 -33678 -10620
rect -33660 -10602 -33624 -10593
rect -33660 -10620 -33651 -10602
rect -33633 -10620 -33624 -10602
rect -33426 -10611 -33381 -10584
rect -33363 -10566 -33309 -10557
rect -33363 -10593 -33345 -10566
rect -33318 -10593 -33309 -10566
rect -33363 -10611 -33309 -10593
rect -33660 -10638 -33624 -10620
rect -35424 -11511 -35415 -11484
rect -35388 -11511 -35379 -11484
rect -35874 -11529 -35838 -11520
rect -35874 -11547 -35865 -11529
rect -35847 -11547 -35838 -11529
rect -35874 -11565 -35838 -11547
rect -35820 -11538 -35757 -11520
rect -35820 -11556 -35811 -11538
rect -35793 -11556 -35757 -11538
rect -35820 -11565 -35757 -11556
rect -35721 -11529 -35676 -11520
rect -35721 -11547 -35712 -11529
rect -35694 -11547 -35676 -11529
rect -35721 -11565 -35676 -11547
rect -35658 -11529 -35622 -11520
rect -35658 -11547 -35649 -11529
rect -35631 -11547 -35622 -11529
rect -35424 -11538 -35379 -11511
rect -35361 -11493 -35307 -11484
rect -35361 -11520 -35343 -11493
rect -35316 -11520 -35307 -11493
rect -35361 -11538 -35307 -11520
rect -35658 -11565 -35622 -11547
rect -35424 -11979 -35415 -11952
rect -35388 -11979 -35379 -11952
rect -35874 -11997 -35838 -11988
rect -35874 -12015 -35865 -11997
rect -35847 -12015 -35838 -11997
rect -35874 -12033 -35838 -12015
rect -35820 -12006 -35757 -11988
rect -35820 -12024 -35811 -12006
rect -35793 -12024 -35757 -12006
rect -35820 -12033 -35757 -12024
rect -35721 -11997 -35676 -11988
rect -35721 -12015 -35712 -11997
rect -35694 -12015 -35676 -11997
rect -35721 -12033 -35676 -12015
rect -35658 -11997 -35622 -11988
rect -35658 -12015 -35649 -11997
rect -35631 -12015 -35622 -11997
rect -35424 -12006 -35379 -11979
rect -35361 -11961 -35307 -11952
rect -35361 -11988 -35343 -11961
rect -35316 -11988 -35307 -11961
rect -35361 -12006 -35307 -11988
rect -35658 -12033 -35622 -12015
rect -33426 -10998 -33417 -10971
rect -33390 -10998 -33381 -10971
rect -33876 -11016 -33840 -11007
rect -33876 -11034 -33867 -11016
rect -33849 -11034 -33840 -11016
rect -33876 -11052 -33840 -11034
rect -33822 -11025 -33759 -11007
rect -33822 -11043 -33813 -11025
rect -33795 -11043 -33759 -11025
rect -33822 -11052 -33759 -11043
rect -33723 -11016 -33678 -11007
rect -33723 -11034 -33714 -11016
rect -33696 -11034 -33678 -11016
rect -33723 -11052 -33678 -11034
rect -33660 -11016 -33624 -11007
rect -33660 -11034 -33651 -11016
rect -33633 -11034 -33624 -11016
rect -33426 -11025 -33381 -10998
rect -33363 -10980 -33309 -10971
rect -33363 -11007 -33345 -10980
rect -33318 -11007 -33309 -10980
rect -33363 -11025 -33309 -11007
rect -33660 -11052 -33624 -11034
rect -29871 -7092 -29808 -7083
rect -29871 -7128 -29862 -7092
rect -29826 -7128 -29808 -7092
rect -29871 -7137 -29808 -7128
rect -29871 -7164 -29808 -7155
rect -29871 -7200 -29862 -7164
rect -29826 -7200 -29808 -7164
rect -29871 -7209 -29808 -7200
rect -29871 -7263 -29808 -7254
rect -29871 -7299 -29862 -7263
rect -29826 -7299 -29808 -7263
rect -29871 -7308 -29808 -7299
rect -29520 -7218 -29511 -7191
rect -29484 -7218 -29475 -7191
rect -29520 -7245 -29475 -7218
rect -29457 -7200 -29403 -7191
rect -29457 -7227 -29439 -7200
rect -29412 -7227 -29403 -7200
rect -29457 -7245 -29403 -7227
rect -29871 -7335 -29808 -7326
rect -29871 -7371 -29862 -7335
rect -29826 -7371 -29808 -7335
rect -29871 -7380 -29808 -7371
rect -29871 -7452 -29808 -7443
rect -29871 -7488 -29862 -7452
rect -29826 -7488 -29808 -7452
rect -29871 -7506 -29808 -7488
rect -29871 -7533 -29808 -7524
rect -29871 -7569 -29862 -7533
rect -29826 -7569 -29808 -7533
rect -29871 -7578 -29808 -7569
rect -29871 -7614 -29808 -7605
rect -29871 -7650 -29862 -7614
rect -29826 -7650 -29808 -7614
rect -29871 -7668 -29808 -7650
rect -29871 -7695 -29808 -7686
rect -29871 -7731 -29862 -7695
rect -29826 -7731 -29808 -7695
rect -29871 -7740 -29808 -7731
rect -29871 -8631 -29808 -8622
rect -29871 -8667 -29862 -8631
rect -29826 -8667 -29808 -8631
rect -29871 -8676 -29808 -8667
rect -29871 -8703 -29808 -8694
rect -29871 -8739 -29862 -8703
rect -29826 -8739 -29808 -8703
rect -29871 -8748 -29808 -8739
rect -29871 -8802 -29808 -8793
rect -29871 -8838 -29862 -8802
rect -29826 -8838 -29808 -8802
rect -29871 -8847 -29808 -8838
rect -28836 -7128 -28791 -7119
rect -28836 -7155 -28827 -7128
rect -28800 -7155 -28791 -7128
rect -28836 -7173 -28791 -7155
rect -28773 -7137 -28728 -7119
rect -28773 -7164 -28764 -7137
rect -28737 -7164 -28728 -7137
rect -28773 -7173 -28728 -7164
rect -28710 -7128 -28665 -7119
rect -28710 -7155 -28701 -7128
rect -28674 -7155 -28665 -7128
rect -28710 -7173 -28665 -7155
rect -28647 -7137 -28593 -7119
rect -28647 -7164 -28638 -7137
rect -28611 -7164 -28593 -7137
rect -28647 -7173 -28593 -7164
rect -28575 -7128 -28521 -7119
rect -28575 -7155 -28557 -7128
rect -28530 -7155 -28521 -7128
rect -28575 -7173 -28521 -7155
rect -28503 -7137 -28458 -7119
rect -28503 -7164 -28494 -7137
rect -28467 -7164 -28458 -7137
rect -28503 -7173 -28458 -7164
rect -28440 -7128 -28395 -7119
rect -28440 -7155 -28431 -7128
rect -28404 -7155 -28395 -7128
rect -28440 -7173 -28395 -7155
rect -28377 -7137 -28332 -7119
rect -28377 -7164 -28368 -7137
rect -28341 -7164 -28332 -7137
rect -28377 -7173 -28332 -7164
rect -28314 -7128 -28260 -7119
rect -28314 -7155 -28305 -7128
rect -28278 -7155 -28260 -7128
rect -28314 -7173 -28260 -7155
rect -28242 -7137 -28107 -7119
rect -28242 -7164 -28233 -7137
rect -28206 -7164 -28107 -7137
rect -28242 -7173 -28107 -7164
rect -28053 -7146 -28035 -7119
rect -28008 -7146 -27999 -7119
rect -28053 -7173 -27999 -7146
rect -27981 -7137 -27936 -7119
rect -27981 -7164 -27972 -7137
rect -27945 -7164 -27936 -7137
rect -27981 -7173 -27936 -7164
rect -29241 -7218 -29232 -7191
rect -29205 -7218 -29196 -7191
rect -29241 -7245 -29196 -7218
rect -29178 -7200 -29124 -7191
rect -29178 -7227 -29160 -7200
rect -29133 -7227 -29124 -7200
rect -29178 -7245 -29124 -7227
rect -29520 -8757 -29511 -8730
rect -29484 -8757 -29475 -8730
rect -29520 -8784 -29475 -8757
rect -29457 -8739 -29403 -8730
rect -29457 -8766 -29439 -8739
rect -29412 -8766 -29403 -8739
rect -29457 -8784 -29403 -8766
rect -29871 -8874 -29808 -8865
rect -29871 -8910 -29862 -8874
rect -29826 -8910 -29808 -8874
rect -29871 -8919 -29808 -8910
rect -29871 -8991 -29808 -8982
rect -29871 -9027 -29862 -8991
rect -29826 -9027 -29808 -8991
rect -29871 -9045 -29808 -9027
rect -29871 -9072 -29808 -9063
rect -29871 -9108 -29862 -9072
rect -29826 -9108 -29808 -9072
rect -29871 -9117 -29808 -9108
rect -29871 -9153 -29808 -9144
rect -29871 -9189 -29862 -9153
rect -29826 -9189 -29808 -9153
rect -29871 -9207 -29808 -9189
rect -29871 -9234 -29808 -9225
rect -29871 -9270 -29862 -9234
rect -29826 -9270 -29808 -9234
rect -29871 -9279 -29808 -9270
rect -29871 -9576 -29808 -9567
rect -29871 -9612 -29862 -9576
rect -29826 -9612 -29808 -9576
rect -29871 -9621 -29808 -9612
rect -29871 -9648 -29808 -9639
rect -29871 -9684 -29862 -9648
rect -29826 -9684 -29808 -9648
rect -29871 -9693 -29808 -9684
rect -29871 -9747 -29808 -9738
rect -29871 -9783 -29862 -9747
rect -29826 -9783 -29808 -9747
rect -29871 -9792 -29808 -9783
rect -29520 -9702 -29511 -9675
rect -29484 -9702 -29475 -9675
rect -29520 -9729 -29475 -9702
rect -29457 -9684 -29403 -9675
rect -29457 -9711 -29439 -9684
rect -29412 -9711 -29403 -9684
rect -29457 -9729 -29403 -9711
rect -29871 -9819 -29808 -9810
rect -29871 -9855 -29862 -9819
rect -29826 -9855 -29808 -9819
rect -29871 -9864 -29808 -9855
rect -29871 -9936 -29808 -9927
rect -29871 -9972 -29862 -9936
rect -29826 -9972 -29808 -9936
rect -29871 -9990 -29808 -9972
rect -29871 -10017 -29808 -10008
rect -29871 -10053 -29862 -10017
rect -29826 -10053 -29808 -10017
rect -29871 -10062 -29808 -10053
rect -29871 -10098 -29808 -10089
rect -29871 -10134 -29862 -10098
rect -29826 -10134 -29808 -10098
rect -26415 -9765 -26406 -9738
rect -26379 -9765 -26370 -9738
rect -28215 -9783 -28170 -9774
rect -28215 -9810 -28206 -9783
rect -28179 -9810 -28170 -9783
rect -28215 -9828 -28170 -9810
rect -28152 -9792 -28107 -9774
rect -28152 -9819 -28143 -9792
rect -28116 -9819 -28107 -9792
rect -28152 -9828 -28107 -9819
rect -28089 -9783 -28044 -9774
rect -28089 -9810 -28080 -9783
rect -28053 -9810 -28044 -9783
rect -28089 -9828 -28044 -9810
rect -28026 -9792 -27972 -9774
rect -28026 -9819 -28017 -9792
rect -27990 -9819 -27972 -9792
rect -28026 -9828 -27972 -9819
rect -27954 -9783 -27900 -9774
rect -27954 -9810 -27936 -9783
rect -27909 -9810 -27900 -9783
rect -27954 -9828 -27900 -9810
rect -27882 -9792 -27837 -9774
rect -27882 -9819 -27873 -9792
rect -27846 -9819 -27837 -9792
rect -27882 -9828 -27837 -9819
rect -27819 -9783 -27774 -9774
rect -27819 -9810 -27810 -9783
rect -27783 -9810 -27774 -9783
rect -27819 -9828 -27774 -9810
rect -27756 -9792 -27711 -9774
rect -27756 -9819 -27747 -9792
rect -27720 -9819 -27711 -9792
rect -27756 -9828 -27711 -9819
rect -27693 -9783 -27639 -9774
rect -27693 -9810 -27684 -9783
rect -27657 -9810 -27639 -9783
rect -27693 -9828 -27639 -9810
rect -27621 -9792 -27486 -9774
rect -27621 -9819 -27612 -9792
rect -27585 -9819 -27486 -9792
rect -27621 -9828 -27486 -9819
rect -27432 -9801 -27414 -9774
rect -27387 -9801 -27378 -9774
rect -27432 -9828 -27378 -9801
rect -27360 -9792 -27315 -9774
rect -27360 -9819 -27351 -9792
rect -27324 -9819 -27315 -9792
rect -26865 -9783 -26829 -9774
rect -26865 -9801 -26856 -9783
rect -26838 -9801 -26829 -9783
rect -26865 -9819 -26829 -9801
rect -26811 -9792 -26748 -9774
rect -26811 -9810 -26802 -9792
rect -26784 -9810 -26748 -9792
rect -26811 -9819 -26748 -9810
rect -26712 -9783 -26667 -9774
rect -26712 -9801 -26703 -9783
rect -26685 -9801 -26667 -9783
rect -26712 -9819 -26667 -9801
rect -26649 -9783 -26613 -9774
rect -26649 -9801 -26640 -9783
rect -26622 -9801 -26613 -9783
rect -26415 -9792 -26370 -9765
rect -26352 -9747 -26298 -9738
rect -26352 -9774 -26334 -9747
rect -26307 -9774 -26298 -9747
rect -26352 -9792 -26298 -9774
rect -26649 -9819 -26613 -9801
rect -27360 -9828 -27315 -9819
rect -29871 -10152 -29808 -10134
rect -29871 -10179 -29808 -10170
rect -29871 -10215 -29862 -10179
rect -29826 -10215 -29808 -10179
rect -29871 -10224 -29808 -10215
rect -29871 -10593 -29808 -10584
rect -29871 -10629 -29862 -10593
rect -29826 -10629 -29808 -10593
rect -29871 -10638 -29808 -10629
rect -29871 -10665 -29808 -10656
rect -29871 -10701 -29862 -10665
rect -29826 -10701 -29808 -10665
rect -29871 -10710 -29808 -10701
rect -29871 -10764 -29808 -10755
rect -29871 -10800 -29862 -10764
rect -29826 -10800 -29808 -10764
rect -29871 -10809 -29808 -10800
rect -29520 -10719 -29511 -10692
rect -29484 -10719 -29475 -10692
rect -29520 -10746 -29475 -10719
rect -29457 -10701 -29403 -10692
rect -29457 -10728 -29439 -10701
rect -29412 -10728 -29403 -10701
rect -29457 -10746 -29403 -10728
rect -29871 -10836 -29808 -10827
rect -29871 -10872 -29862 -10836
rect -29826 -10872 -29808 -10836
rect -29871 -10881 -29808 -10872
rect -29871 -10953 -29808 -10944
rect -29871 -10989 -29862 -10953
rect -29826 -10989 -29808 -10953
rect -29871 -11007 -29808 -10989
rect -29871 -11034 -29808 -11025
rect -29871 -11070 -29862 -11034
rect -29826 -11070 -29808 -11034
rect -29871 -11079 -29808 -11070
rect -29871 -11115 -29808 -11106
rect -29871 -11151 -29862 -11115
rect -29826 -11151 -29808 -11115
rect -29871 -11169 -29808 -11151
rect -29871 -11196 -29808 -11187
rect -29871 -11232 -29862 -11196
rect -29826 -11232 -29808 -11196
rect -29871 -11241 -29808 -11232
rect -33426 -11529 -33417 -11502
rect -33390 -11529 -33381 -11502
rect -33876 -11547 -33840 -11538
rect -33876 -11565 -33867 -11547
rect -33849 -11565 -33840 -11547
rect -33876 -11583 -33840 -11565
rect -33822 -11556 -33759 -11538
rect -33822 -11574 -33813 -11556
rect -33795 -11574 -33759 -11556
rect -33822 -11583 -33759 -11574
rect -33723 -11547 -33678 -11538
rect -33723 -11565 -33714 -11547
rect -33696 -11565 -33678 -11547
rect -33723 -11583 -33678 -11565
rect -33660 -11547 -33624 -11538
rect -33660 -11565 -33651 -11547
rect -33633 -11565 -33624 -11547
rect -33426 -11556 -33381 -11529
rect -33363 -11511 -33309 -11502
rect -33363 -11538 -33345 -11511
rect -33318 -11538 -33309 -11511
rect -33363 -11556 -33309 -11538
rect -33660 -11583 -33624 -11565
rect -36216 -12168 -36207 -12141
rect -36180 -12168 -36171 -12141
rect -36216 -12195 -36171 -12168
rect -36153 -12150 -36099 -12141
rect -36153 -12177 -36135 -12150
rect -36108 -12177 -36099 -12150
rect -36153 -12195 -36099 -12177
rect -35424 -12420 -35415 -12393
rect -35388 -12420 -35379 -12393
rect -35874 -12438 -35838 -12429
rect -35874 -12456 -35865 -12438
rect -35847 -12456 -35838 -12438
rect -36207 -12492 -36198 -12465
rect -36171 -12492 -36162 -12465
rect -36207 -12519 -36162 -12492
rect -36144 -12474 -36090 -12465
rect -35874 -12474 -35838 -12456
rect -35820 -12447 -35757 -12429
rect -35820 -12465 -35811 -12447
rect -35793 -12465 -35757 -12447
rect -35820 -12474 -35757 -12465
rect -35721 -12438 -35676 -12429
rect -35721 -12456 -35712 -12438
rect -35694 -12456 -35676 -12438
rect -35721 -12474 -35676 -12456
rect -35658 -12438 -35622 -12429
rect -35658 -12456 -35649 -12438
rect -35631 -12456 -35622 -12438
rect -35424 -12447 -35379 -12420
rect -35361 -12402 -35307 -12393
rect -35361 -12429 -35343 -12402
rect -35316 -12429 -35307 -12402
rect -29871 -11889 -29808 -11880
rect -29871 -11925 -29862 -11889
rect -29826 -11925 -29808 -11889
rect -29871 -11934 -29808 -11925
rect -33426 -12393 -33417 -12366
rect -33390 -12393 -33381 -12366
rect -35361 -12447 -35307 -12429
rect -33876 -12411 -33840 -12402
rect -33876 -12429 -33867 -12411
rect -33849 -12429 -33840 -12411
rect -35658 -12474 -35622 -12456
rect -36144 -12501 -36126 -12474
rect -36099 -12501 -36090 -12474
rect -36144 -12519 -36090 -12501
rect -33876 -12447 -33840 -12429
rect -33822 -12420 -33759 -12402
rect -33822 -12438 -33813 -12420
rect -33795 -12438 -33759 -12420
rect -33822 -12447 -33759 -12438
rect -33723 -12411 -33678 -12402
rect -33723 -12429 -33714 -12411
rect -33696 -12429 -33678 -12411
rect -33723 -12447 -33678 -12429
rect -33660 -12411 -33624 -12402
rect -33660 -12429 -33651 -12411
rect -33633 -12429 -33624 -12411
rect -33426 -12420 -33381 -12393
rect -33363 -12375 -33309 -12366
rect -33363 -12402 -33345 -12375
rect -33318 -12402 -33309 -12375
rect -33363 -12420 -33309 -12402
rect -33660 -12447 -33624 -12429
rect -35424 -12834 -35415 -12807
rect -35388 -12834 -35379 -12807
rect -35874 -12852 -35838 -12843
rect -35874 -12870 -35865 -12852
rect -35847 -12870 -35838 -12852
rect -35874 -12888 -35838 -12870
rect -35820 -12861 -35757 -12843
rect -35820 -12879 -35811 -12861
rect -35793 -12879 -35757 -12861
rect -35820 -12888 -35757 -12879
rect -35721 -12852 -35676 -12843
rect -35721 -12870 -35712 -12852
rect -35694 -12870 -35676 -12852
rect -35721 -12888 -35676 -12870
rect -35658 -12852 -35622 -12843
rect -35658 -12870 -35649 -12852
rect -35631 -12870 -35622 -12852
rect -35424 -12861 -35379 -12834
rect -35361 -12816 -35307 -12807
rect -35361 -12843 -35343 -12816
rect -35316 -12843 -35307 -12816
rect -35361 -12861 -35307 -12843
rect -35658 -12888 -35622 -12870
rect -29871 -11961 -29808 -11952
rect -29871 -11997 -29862 -11961
rect -29826 -11997 -29808 -11961
rect -29871 -12006 -29808 -11997
rect -29871 -12060 -29808 -12051
rect -29871 -12096 -29862 -12060
rect -29826 -12096 -29808 -12060
rect -29871 -12105 -29808 -12096
rect -29520 -12015 -29511 -11988
rect -29484 -12015 -29475 -11988
rect -29520 -12042 -29475 -12015
rect -29457 -11997 -29403 -11988
rect -29457 -12024 -29439 -11997
rect -29412 -12024 -29403 -11997
rect -29457 -12042 -29403 -12024
rect -29871 -12132 -29808 -12123
rect -29871 -12168 -29862 -12132
rect -29826 -12168 -29808 -12132
rect -29871 -12177 -29808 -12168
rect -29871 -12249 -29808 -12240
rect -29871 -12285 -29862 -12249
rect -29826 -12285 -29808 -12249
rect -29871 -12303 -29808 -12285
rect -29871 -12330 -29808 -12321
rect -29871 -12366 -29862 -12330
rect -29826 -12366 -29808 -12330
rect -29871 -12375 -29808 -12366
rect -29871 -12411 -29808 -12402
rect -29871 -12447 -29862 -12411
rect -29826 -12447 -29808 -12411
rect -29871 -12465 -29808 -12447
rect -29871 -12492 -29808 -12483
rect -29871 -12528 -29862 -12492
rect -29826 -12528 -29808 -12492
rect -29871 -12537 -29808 -12528
rect -33426 -12888 -33417 -12861
rect -33390 -12888 -33381 -12861
rect -33876 -12906 -33840 -12897
rect -33876 -12924 -33867 -12906
rect -33849 -12924 -33840 -12906
rect -33876 -12942 -33840 -12924
rect -33822 -12915 -33759 -12897
rect -33822 -12933 -33813 -12915
rect -33795 -12933 -33759 -12915
rect -33822 -12942 -33759 -12933
rect -33723 -12906 -33678 -12897
rect -33723 -12924 -33714 -12906
rect -33696 -12924 -33678 -12906
rect -33723 -12942 -33678 -12924
rect -33660 -12906 -33624 -12897
rect -33660 -12924 -33651 -12906
rect -33633 -12924 -33624 -12906
rect -33426 -12915 -33381 -12888
rect -33363 -12870 -33309 -12861
rect -33363 -12897 -33345 -12870
rect -33318 -12897 -33309 -12870
rect -33363 -12915 -33309 -12897
rect -33660 -12942 -33624 -12924
rect -33426 -13302 -33417 -13275
rect -33390 -13302 -33381 -13275
rect -33876 -13320 -33840 -13311
rect -33876 -13338 -33867 -13320
rect -33849 -13338 -33840 -13320
rect -33876 -13356 -33840 -13338
rect -33822 -13329 -33759 -13311
rect -33822 -13347 -33813 -13329
rect -33795 -13347 -33759 -13329
rect -33822 -13356 -33759 -13347
rect -33723 -13320 -33678 -13311
rect -33723 -13338 -33714 -13320
rect -33696 -13338 -33678 -13320
rect -33723 -13356 -33678 -13338
rect -33660 -13320 -33624 -13311
rect -33660 -13338 -33651 -13320
rect -33633 -13338 -33624 -13320
rect -33426 -13329 -33381 -13302
rect -33363 -13284 -33309 -13275
rect -33363 -13311 -33345 -13284
rect -33318 -13311 -33309 -13284
rect -33363 -13329 -33309 -13311
rect -33660 -13356 -33624 -13338
rect -33426 -13833 -33417 -13806
rect -33390 -13833 -33381 -13806
rect -33876 -13851 -33840 -13842
rect -33876 -13869 -33867 -13851
rect -33849 -13869 -33840 -13851
rect -33876 -13887 -33840 -13869
rect -33822 -13860 -33759 -13842
rect -33822 -13878 -33813 -13860
rect -33795 -13878 -33759 -13860
rect -33822 -13887 -33759 -13878
rect -33723 -13851 -33678 -13842
rect -33723 -13869 -33714 -13851
rect -33696 -13869 -33678 -13851
rect -33723 -13887 -33678 -13869
rect -33660 -13851 -33624 -13842
rect -33660 -13869 -33651 -13851
rect -33633 -13869 -33624 -13851
rect -33426 -13860 -33381 -13833
rect -33363 -13815 -33309 -13806
rect -33363 -13842 -33345 -13815
rect -33318 -13842 -33309 -13815
rect -33363 -13860 -33309 -13842
rect -31455 -13842 -31446 -13815
rect -31419 -13842 -31410 -13815
rect -31905 -13860 -31869 -13851
rect -33660 -13887 -33624 -13869
rect -31905 -13878 -31896 -13860
rect -31878 -13878 -31869 -13860
rect -31905 -13896 -31869 -13878
rect -31851 -13869 -31788 -13851
rect -31851 -13887 -31842 -13869
rect -31824 -13887 -31788 -13869
rect -31851 -13896 -31788 -13887
rect -31752 -13860 -31707 -13851
rect -31752 -13878 -31743 -13860
rect -31725 -13878 -31707 -13860
rect -31752 -13896 -31707 -13878
rect -31689 -13860 -31653 -13851
rect -31689 -13878 -31680 -13860
rect -31662 -13878 -31653 -13860
rect -31455 -13869 -31410 -13842
rect -31392 -13824 -31338 -13815
rect -31392 -13851 -31374 -13824
rect -31347 -13851 -31338 -13824
rect -31392 -13869 -31338 -13851
rect -31689 -13896 -31653 -13878
rect -33426 -14328 -33417 -14301
rect -33390 -14328 -33381 -14301
rect -33876 -14346 -33840 -14337
rect -33876 -14364 -33867 -14346
rect -33849 -14364 -33840 -14346
rect -33876 -14382 -33840 -14364
rect -33822 -14355 -33759 -14337
rect -33822 -14373 -33813 -14355
rect -33795 -14373 -33759 -14355
rect -33822 -14382 -33759 -14373
rect -33723 -14346 -33678 -14337
rect -33723 -14364 -33714 -14346
rect -33696 -14364 -33678 -14346
rect -33723 -14382 -33678 -14364
rect -33660 -14346 -33624 -14337
rect -33660 -14364 -33651 -14346
rect -33633 -14364 -33624 -14346
rect -33426 -14355 -33381 -14328
rect -33363 -14310 -33309 -14301
rect -33363 -14337 -33345 -14310
rect -33318 -14337 -33309 -14310
rect -31455 -14319 -31446 -14292
rect -31419 -14319 -31410 -14292
rect -33363 -14355 -33309 -14337
rect -31905 -14337 -31869 -14328
rect -31905 -14355 -31896 -14337
rect -31878 -14355 -31869 -14337
rect -33660 -14382 -33624 -14364
rect -31905 -14373 -31869 -14355
rect -31851 -14346 -31788 -14328
rect -31851 -14364 -31842 -14346
rect -31824 -14364 -31788 -14346
rect -31851 -14373 -31788 -14364
rect -31752 -14337 -31707 -14328
rect -31752 -14355 -31743 -14337
rect -31725 -14355 -31707 -14337
rect -31752 -14373 -31707 -14355
rect -31689 -14337 -31653 -14328
rect -31689 -14355 -31680 -14337
rect -31662 -14355 -31653 -14337
rect -31455 -14346 -31410 -14319
rect -31392 -14301 -31338 -14292
rect -31392 -14328 -31374 -14301
rect -31347 -14328 -31338 -14301
rect -31392 -14346 -31338 -14328
rect -31689 -14373 -31653 -14355
rect -31455 -14715 -31446 -14688
rect -31419 -14715 -31410 -14688
rect -31905 -14733 -31869 -14724
rect -31905 -14751 -31896 -14733
rect -31878 -14751 -31869 -14733
rect -31905 -14769 -31869 -14751
rect -31851 -14742 -31788 -14724
rect -31851 -14760 -31842 -14742
rect -31824 -14760 -31788 -14742
rect -31851 -14769 -31788 -14760
rect -31752 -14733 -31707 -14724
rect -31752 -14751 -31743 -14733
rect -31725 -14751 -31707 -14733
rect -31752 -14769 -31707 -14751
rect -31689 -14733 -31653 -14724
rect -31689 -14751 -31680 -14733
rect -31662 -14751 -31653 -14733
rect -31455 -14742 -31410 -14715
rect -31392 -14697 -31338 -14688
rect -31392 -14724 -31374 -14697
rect -31347 -14724 -31338 -14697
rect -31392 -14742 -31338 -14724
rect -31689 -14769 -31653 -14751
rect -33426 -14823 -33417 -14796
rect -33390 -14823 -33381 -14796
rect -33876 -14841 -33840 -14832
rect -33876 -14859 -33867 -14841
rect -33849 -14859 -33840 -14841
rect -33876 -14877 -33840 -14859
rect -33822 -14850 -33759 -14832
rect -33822 -14868 -33813 -14850
rect -33795 -14868 -33759 -14850
rect -33822 -14877 -33759 -14868
rect -33723 -14841 -33678 -14832
rect -33723 -14859 -33714 -14841
rect -33696 -14859 -33678 -14841
rect -33723 -14877 -33678 -14859
rect -33660 -14841 -33624 -14832
rect -33660 -14859 -33651 -14841
rect -33633 -14859 -33624 -14841
rect -33426 -14850 -33381 -14823
rect -33363 -14805 -33309 -14796
rect -33363 -14832 -33345 -14805
rect -33318 -14832 -33309 -14805
rect -33363 -14850 -33309 -14832
rect -33660 -14877 -33624 -14859
rect -31455 -15183 -31446 -15156
rect -31419 -15183 -31410 -15156
rect -31905 -15201 -31869 -15192
rect -33426 -15237 -33417 -15210
rect -33390 -15237 -33381 -15210
rect -33876 -15255 -33840 -15246
rect -33876 -15273 -33867 -15255
rect -33849 -15273 -33840 -15255
rect -33876 -15291 -33840 -15273
rect -33822 -15264 -33759 -15246
rect -33822 -15282 -33813 -15264
rect -33795 -15282 -33759 -15264
rect -33822 -15291 -33759 -15282
rect -33723 -15255 -33678 -15246
rect -33723 -15273 -33714 -15255
rect -33696 -15273 -33678 -15255
rect -33723 -15291 -33678 -15273
rect -33660 -15255 -33624 -15246
rect -33660 -15273 -33651 -15255
rect -33633 -15273 -33624 -15255
rect -33426 -15264 -33381 -15237
rect -33363 -15219 -33309 -15210
rect -33363 -15246 -33345 -15219
rect -33318 -15246 -33309 -15219
rect -31905 -15219 -31896 -15201
rect -31878 -15219 -31869 -15201
rect -31905 -15237 -31869 -15219
rect -31851 -15210 -31788 -15192
rect -31851 -15228 -31842 -15210
rect -31824 -15228 -31788 -15210
rect -31851 -15237 -31788 -15228
rect -31752 -15201 -31707 -15192
rect -31752 -15219 -31743 -15201
rect -31725 -15219 -31707 -15201
rect -31752 -15237 -31707 -15219
rect -31689 -15201 -31653 -15192
rect -31689 -15219 -31680 -15201
rect -31662 -15219 -31653 -15201
rect -31455 -15210 -31410 -15183
rect -31392 -15165 -31338 -15156
rect -31392 -15192 -31374 -15165
rect -31347 -15192 -31338 -15165
rect -31392 -15210 -31338 -15192
rect -31689 -15237 -31653 -15219
rect -33363 -15264 -33309 -15246
rect -33660 -15291 -33624 -15273
rect -33426 -15768 -33417 -15741
rect -33390 -15768 -33381 -15741
rect -33876 -15786 -33840 -15777
rect -33876 -15804 -33867 -15786
rect -33849 -15804 -33840 -15786
rect -33876 -15822 -33840 -15804
rect -33822 -15795 -33759 -15777
rect -33822 -15813 -33813 -15795
rect -33795 -15813 -33759 -15795
rect -33822 -15822 -33759 -15813
rect -33723 -15786 -33678 -15777
rect -33723 -15804 -33714 -15786
rect -33696 -15804 -33678 -15786
rect -33723 -15822 -33678 -15804
rect -33660 -15786 -33624 -15777
rect -33660 -15804 -33651 -15786
rect -33633 -15804 -33624 -15786
rect -33426 -15795 -33381 -15768
rect -33363 -15750 -33309 -15741
rect -33363 -15777 -33345 -15750
rect -33318 -15777 -33309 -15750
rect -33363 -15795 -33309 -15777
rect -33660 -15822 -33624 -15804
<< ndcontact >>
rect -30474 10296 -30438 10332
rect -30474 10224 -30438 10260
rect -30474 10125 -30438 10161
rect -29664 10296 -29628 10332
rect -30474 10053 -30438 10089
rect -30474 9936 -30438 9972
rect -30474 9855 -30438 9891
rect -30474 9774 -30438 9810
rect -30474 9693 -30438 9729
rect -29664 10224 -29628 10260
rect -29664 10125 -29628 10161
rect -28782 10296 -28746 10332
rect -29664 10053 -29628 10089
rect -29664 9936 -29628 9972
rect -29664 9855 -29628 9891
rect -29664 9774 -29628 9810
rect -29664 9693 -29628 9729
rect -28782 10224 -28746 10260
rect -28782 10125 -28746 10161
rect -28782 10053 -28746 10089
rect -28782 9936 -28746 9972
rect -28782 9855 -28746 9891
rect -28782 9774 -28746 9810
rect -28782 9693 -28746 9729
rect -29907 9216 -29880 9243
rect -29835 9225 -29808 9252
rect -30357 9171 -30339 9189
rect -30141 9180 -30123 9198
rect -29331 9234 -29313 9252
rect -29115 9243 -29097 9261
rect -28881 9279 -28854 9306
rect -28809 9288 -28782 9315
rect -29682 8829 -29664 8847
rect -29628 8829 -29610 8847
rect -29592 8829 -29574 8847
rect -29538 8829 -29520 8847
rect -29466 8829 -29448 8847
rect -29412 8829 -29394 8847
rect -30474 8199 -30438 8235
rect -30474 8127 -30438 8163
rect -30474 8028 -30438 8064
rect -29664 8199 -29628 8235
rect -30474 7956 -30438 7992
rect -30474 7839 -30438 7875
rect -30474 7758 -30438 7794
rect -30474 7677 -30438 7713
rect -30474 7596 -30438 7632
rect -29664 8127 -29628 8163
rect -29664 8028 -29628 8064
rect -28782 8199 -28746 8235
rect -29664 7956 -29628 7992
rect -29664 7839 -29628 7875
rect -29664 7758 -29628 7794
rect -29664 7677 -29628 7713
rect -29664 7596 -29628 7632
rect -28782 8127 -28746 8163
rect -28782 8028 -28746 8064
rect -28782 7956 -28746 7992
rect -28782 7839 -28746 7875
rect -28782 7758 -28746 7794
rect -28782 7677 -28746 7713
rect -28782 7596 -28746 7632
rect -29907 7119 -29880 7146
rect -29835 7128 -29808 7155
rect -30357 7074 -30339 7092
rect -30141 7083 -30123 7101
rect -29331 7137 -29313 7155
rect -29115 7146 -29097 7164
rect -28881 7182 -28854 7209
rect -28809 7191 -28782 7218
rect -29682 6732 -29664 6750
rect -29628 6732 -29610 6750
rect -29592 6732 -29574 6750
rect -29538 6732 -29520 6750
rect -29466 6732 -29448 6750
rect -29412 6732 -29394 6750
rect -30474 6084 -30438 6120
rect -30474 6012 -30438 6048
rect -30474 5913 -30438 5949
rect -29664 6084 -29628 6120
rect -30474 5841 -30438 5877
rect -30474 5724 -30438 5760
rect -30474 5643 -30438 5679
rect -30474 5562 -30438 5598
rect -30474 5481 -30438 5517
rect -29664 6012 -29628 6048
rect -29664 5913 -29628 5949
rect -28782 6084 -28746 6120
rect -29664 5841 -29628 5877
rect -29664 5724 -29628 5760
rect -29664 5643 -29628 5679
rect -29664 5562 -29628 5598
rect -29664 5481 -29628 5517
rect -28782 6012 -28746 6048
rect -28782 5913 -28746 5949
rect -28782 5841 -28746 5877
rect -28782 5724 -28746 5760
rect -28782 5643 -28746 5679
rect -28782 5562 -28746 5598
rect -28782 5481 -28746 5517
rect -29907 5004 -29880 5031
rect -29835 5013 -29808 5040
rect -30357 4959 -30339 4977
rect -30141 4968 -30123 4986
rect -29331 5022 -29313 5040
rect -29115 5031 -29097 5049
rect -28881 5067 -28854 5094
rect -28809 5076 -28782 5103
rect -29682 4617 -29664 4635
rect -29628 4617 -29610 4635
rect -29592 4617 -29574 4635
rect -29538 4617 -29520 4635
rect -29466 4617 -29448 4635
rect -29412 4617 -29394 4635
rect -30474 4149 -30438 4185
rect -30474 4077 -30438 4113
rect -30474 3978 -30438 4014
rect -29664 4149 -29628 4185
rect -30474 3906 -30438 3942
rect -30474 3789 -30438 3825
rect -30474 3708 -30438 3744
rect -30474 3627 -30438 3663
rect -30474 3546 -30438 3582
rect -29664 4077 -29628 4113
rect -29664 3978 -29628 4014
rect -28782 4149 -28746 4185
rect -29664 3906 -29628 3942
rect -29664 3789 -29628 3825
rect -29664 3708 -29628 3744
rect -29664 3627 -29628 3663
rect -29664 3546 -29628 3582
rect -28782 4077 -28746 4113
rect -28782 3978 -28746 4014
rect -28782 3906 -28746 3942
rect -28782 3789 -28746 3825
rect -28782 3708 -28746 3744
rect -28782 3627 -28746 3663
rect -28782 3546 -28746 3582
rect -29907 3069 -29880 3096
rect -29835 3078 -29808 3105
rect -30357 3024 -30339 3042
rect -30141 3033 -30123 3051
rect -29331 3087 -29313 3105
rect -29115 3096 -29097 3114
rect -28881 3132 -28854 3159
rect -28809 3141 -28782 3168
rect -29682 2682 -29664 2700
rect -29628 2682 -29610 2700
rect -29592 2682 -29574 2700
rect -29538 2682 -29520 2700
rect -29466 2682 -29448 2700
rect -29412 2682 -29394 2700
rect -30114 459 -30078 495
rect -30114 387 -30078 423
rect -30114 288 -30078 324
rect -30114 216 -30078 252
rect -29511 234 -29484 261
rect -29439 243 -29412 270
rect -30114 99 -30078 135
rect -30114 18 -30078 54
rect -30114 -63 -30078 -27
rect -30114 -144 -30078 -108
rect -29142 -72 -29115 -45
rect -29070 -63 -29043 -36
rect -28305 -36 -28278 -9
rect -28233 -27 -28206 0
rect -28755 -81 -28737 -63
rect -28539 -72 -28521 -54
rect -33435 -450 -33408 -423
rect -33363 -441 -33336 -414
rect -33885 -495 -33867 -477
rect -33669 -486 -33651 -468
rect -30114 -486 -30078 -450
rect -33435 -945 -33408 -918
rect -33363 -936 -33336 -909
rect -33885 -990 -33867 -972
rect -33669 -981 -33651 -963
rect -34452 -1224 -34434 -1206
rect -34398 -1224 -34380 -1206
rect -34362 -1224 -34344 -1206
rect -34308 -1224 -34290 -1206
rect -34236 -1224 -34218 -1206
rect -34182 -1224 -34164 -1206
rect -33435 -1359 -33408 -1332
rect -33363 -1350 -33336 -1323
rect -33885 -1404 -33867 -1386
rect -33669 -1395 -33651 -1377
rect -33435 -1890 -33408 -1863
rect -33363 -1881 -33336 -1854
rect -33885 -1935 -33867 -1917
rect -33669 -1926 -33651 -1908
rect -33435 -2457 -33408 -2430
rect -33363 -2448 -33336 -2421
rect -33885 -2502 -33867 -2484
rect -33669 -2493 -33651 -2475
rect -33435 -2952 -33408 -2925
rect -33363 -2943 -33336 -2916
rect -33885 -2997 -33867 -2979
rect -33669 -2988 -33651 -2970
rect -33435 -3366 -33408 -3339
rect -33363 -3357 -33336 -3330
rect -33885 -3411 -33867 -3393
rect -33669 -3402 -33651 -3384
rect -33435 -3897 -33408 -3870
rect -33363 -3888 -33336 -3861
rect -33885 -3942 -33867 -3924
rect -33669 -3933 -33651 -3915
rect -30114 -558 -30078 -522
rect -30114 -657 -30078 -621
rect -30114 -729 -30078 -693
rect -29511 -711 -29484 -684
rect -29439 -702 -29412 -675
rect -30114 -846 -30078 -810
rect -30114 -927 -30078 -891
rect -29160 -882 -29133 -855
rect -29088 -873 -29061 -846
rect -28377 -846 -28350 -819
rect -28305 -837 -28278 -810
rect -27549 -846 -27522 -819
rect -27477 -837 -27450 -810
rect -28827 -891 -28809 -873
rect -28611 -882 -28593 -864
rect -27999 -891 -27981 -873
rect -27783 -882 -27765 -864
rect -27126 -882 -27108 -864
rect -27063 -882 -27045 -864
rect -27027 -882 -27009 -864
rect -26973 -882 -26955 -864
rect -26937 -882 -26919 -864
rect -26883 -882 -26865 -864
rect -26847 -882 -26829 -864
rect -26793 -882 -26775 -864
rect -26721 -882 -26703 -864
rect -26667 -882 -26649 -864
rect -30114 -1008 -30078 -972
rect -30114 -1089 -30078 -1053
rect -30114 -1503 -30078 -1467
rect -30114 -1575 -30078 -1539
rect -30114 -1674 -30078 -1638
rect -30114 -1746 -30078 -1710
rect -29511 -1728 -29484 -1701
rect -29439 -1719 -29412 -1692
rect -29178 -1728 -29151 -1701
rect -29106 -1719 -29079 -1692
rect -28674 -1701 -28647 -1674
rect -28053 -1701 -28026 -1674
rect -27882 -1701 -27855 -1674
rect -27819 -1701 -27792 -1674
rect -30114 -1863 -30078 -1827
rect -30114 -1944 -30078 -1908
rect -30114 -2025 -30078 -1989
rect -30114 -2106 -30078 -2070
rect -30114 -2799 -30078 -2763
rect -30114 -2871 -30078 -2835
rect -30114 -2970 -30078 -2934
rect -30114 -3042 -30078 -3006
rect -29511 -3024 -29484 -2997
rect -29439 -3015 -29412 -2988
rect -29232 -3024 -29205 -2997
rect -29160 -3015 -29133 -2988
rect -28827 -2997 -28800 -2970
rect -28206 -2997 -28179 -2970
rect -28035 -2997 -28008 -2970
rect -27972 -2997 -27945 -2970
rect -30114 -3159 -30078 -3123
rect -30114 -3240 -30078 -3204
rect -30114 -3321 -30078 -3285
rect -30114 -3402 -30078 -3366
rect -30114 -3870 -30078 -3834
rect -30114 -3942 -30078 -3906
rect -30114 -4041 -30078 -4005
rect -30114 -4113 -30078 -4077
rect -29511 -4095 -29484 -4068
rect -29439 -4086 -29412 -4059
rect -30114 -4230 -30078 -4194
rect -30114 -4311 -30078 -4275
rect -30114 -4392 -30078 -4356
rect -30114 -4473 -30078 -4437
rect -29142 -4401 -29115 -4374
rect -29070 -4392 -29043 -4365
rect -28305 -4365 -28278 -4338
rect -28233 -4356 -28206 -4329
rect -28755 -4410 -28737 -4392
rect -28539 -4401 -28521 -4383
rect -30114 -4815 -30078 -4779
rect -30114 -4887 -30078 -4851
rect -30114 -4986 -30078 -4950
rect -30114 -5058 -30078 -5022
rect -29511 -5040 -29484 -5013
rect -29439 -5031 -29412 -5004
rect -30114 -5175 -30078 -5139
rect -30114 -5256 -30078 -5220
rect -29160 -5211 -29133 -5184
rect -29088 -5202 -29061 -5175
rect -28377 -5175 -28350 -5148
rect -28305 -5166 -28278 -5139
rect -27549 -5175 -27522 -5148
rect -27477 -5166 -27450 -5139
rect -28827 -5220 -28809 -5202
rect -28611 -5211 -28593 -5193
rect -27999 -5220 -27981 -5202
rect -27783 -5211 -27765 -5193
rect -27126 -5211 -27108 -5193
rect -27063 -5211 -27045 -5193
rect -27027 -5211 -27009 -5193
rect -26973 -5211 -26955 -5193
rect -26937 -5211 -26919 -5193
rect -26883 -5211 -26865 -5193
rect -26847 -5211 -26829 -5193
rect -26793 -5211 -26775 -5193
rect -26721 -5211 -26703 -5193
rect -26667 -5211 -26649 -5193
rect -30114 -5337 -30078 -5301
rect -30114 -5418 -30078 -5382
rect -30114 -5832 -30078 -5796
rect -30114 -5904 -30078 -5868
rect -30114 -6003 -30078 -5967
rect -30114 -6075 -30078 -6039
rect -29511 -6057 -29484 -6030
rect -29439 -6048 -29412 -6021
rect -29178 -6057 -29151 -6030
rect -29106 -6048 -29079 -6021
rect -28674 -6030 -28647 -6003
rect -28053 -6030 -28026 -6003
rect -27882 -6030 -27855 -6003
rect -27819 -6030 -27792 -6003
rect -30114 -6192 -30078 -6156
rect -30114 -6273 -30078 -6237
rect -30114 -6354 -30078 -6318
rect -30114 -6435 -30078 -6399
rect -33417 -8307 -33390 -8280
rect -33345 -8298 -33318 -8271
rect -33867 -8352 -33849 -8334
rect -33651 -8343 -33633 -8325
rect -33417 -8802 -33390 -8775
rect -33345 -8793 -33318 -8766
rect -33867 -8847 -33849 -8829
rect -33651 -8838 -33633 -8820
rect -33417 -9216 -33390 -9189
rect -33345 -9207 -33318 -9180
rect -33867 -9261 -33849 -9243
rect -33651 -9252 -33633 -9234
rect -33417 -9747 -33390 -9720
rect -33345 -9738 -33318 -9711
rect -33867 -9792 -33849 -9774
rect -33651 -9783 -33633 -9765
rect -33417 -10224 -33390 -10197
rect -33345 -10215 -33318 -10188
rect -33867 -10269 -33849 -10251
rect -33651 -10260 -33633 -10242
rect -35415 -11646 -35388 -11619
rect -35343 -11637 -35316 -11610
rect -35865 -11691 -35847 -11673
rect -35649 -11682 -35631 -11664
rect -33417 -10719 -33390 -10692
rect -33345 -10710 -33318 -10683
rect -33867 -10764 -33849 -10746
rect -33651 -10755 -33633 -10737
rect -33417 -11133 -33390 -11106
rect -33345 -11124 -33318 -11097
rect -33867 -11178 -33849 -11160
rect -33651 -11169 -33633 -11151
rect -30114 -7128 -30078 -7092
rect -30114 -7200 -30078 -7164
rect -30114 -7299 -30078 -7263
rect -30114 -7371 -30078 -7335
rect -29511 -7353 -29484 -7326
rect -29439 -7344 -29412 -7317
rect -30114 -7488 -30078 -7452
rect -30114 -7569 -30078 -7533
rect -30114 -7650 -30078 -7614
rect -30114 -7731 -30078 -7695
rect -30114 -8667 -30078 -8631
rect -30114 -8739 -30078 -8703
rect -30114 -8838 -30078 -8802
rect -29232 -7353 -29205 -7326
rect -29160 -7344 -29133 -7317
rect -28827 -7326 -28800 -7299
rect -28206 -7326 -28179 -7299
rect -28035 -7326 -28008 -7299
rect -27972 -7326 -27945 -7299
rect -30114 -8910 -30078 -8874
rect -29511 -8892 -29484 -8865
rect -29439 -8883 -29412 -8856
rect -30114 -9027 -30078 -8991
rect -30114 -9108 -30078 -9072
rect -30114 -9189 -30078 -9153
rect -30114 -9270 -30078 -9234
rect -30114 -9612 -30078 -9576
rect -30114 -9684 -30078 -9648
rect -30114 -9783 -30078 -9747
rect -30114 -9855 -30078 -9819
rect -29511 -9837 -29484 -9810
rect -29439 -9828 -29412 -9801
rect -30114 -9972 -30078 -9936
rect -30114 -10053 -30078 -10017
rect -30114 -10134 -30078 -10098
rect -26406 -9900 -26379 -9873
rect -26334 -9891 -26307 -9864
rect -26856 -9945 -26838 -9927
rect -26640 -9936 -26622 -9918
rect -28206 -9981 -28179 -9954
rect -27585 -9981 -27558 -9954
rect -27414 -9981 -27387 -9954
rect -27351 -9981 -27324 -9954
rect -30114 -10215 -30078 -10179
rect -30114 -10629 -30078 -10593
rect -30114 -10701 -30078 -10665
rect -30114 -10800 -30078 -10764
rect -30114 -10872 -30078 -10836
rect -29511 -10854 -29484 -10827
rect -29439 -10845 -29412 -10818
rect -30114 -10989 -30078 -10953
rect -30114 -11070 -30078 -11034
rect -30114 -11151 -30078 -11115
rect -30114 -11232 -30078 -11196
rect -35415 -12114 -35388 -12087
rect -35343 -12105 -35316 -12078
rect -35865 -12159 -35847 -12141
rect -35649 -12150 -35631 -12132
rect -36207 -12303 -36180 -12276
rect -36135 -12294 -36108 -12267
rect -33417 -11664 -33390 -11637
rect -33345 -11655 -33318 -11628
rect -33867 -11709 -33849 -11691
rect -33651 -11700 -33633 -11682
rect -30114 -11925 -30078 -11889
rect -35415 -12555 -35388 -12528
rect -35343 -12546 -35316 -12519
rect -36198 -12627 -36171 -12600
rect -36126 -12618 -36099 -12591
rect -35865 -12600 -35847 -12582
rect -35649 -12591 -35631 -12573
rect -33417 -12528 -33390 -12501
rect -33345 -12519 -33318 -12492
rect -33867 -12573 -33849 -12555
rect -33651 -12564 -33633 -12546
rect -30114 -11997 -30078 -11961
rect -30114 -12096 -30078 -12060
rect -30114 -12168 -30078 -12132
rect -29511 -12150 -29484 -12123
rect -29439 -12141 -29412 -12114
rect -30114 -12285 -30078 -12249
rect -30114 -12366 -30078 -12330
rect -30114 -12447 -30078 -12411
rect -30114 -12528 -30078 -12492
rect -35415 -12969 -35388 -12942
rect -35343 -12960 -35316 -12933
rect -35865 -13014 -35847 -12996
rect -35649 -13005 -35631 -12987
rect -33417 -13023 -33390 -12996
rect -33345 -13014 -33318 -12987
rect -33867 -13068 -33849 -13050
rect -33651 -13059 -33633 -13041
rect -33417 -13437 -33390 -13410
rect -33345 -13428 -33318 -13401
rect -33867 -13482 -33849 -13464
rect -33651 -13473 -33633 -13455
rect -33417 -13968 -33390 -13941
rect -33345 -13959 -33318 -13932
rect -33867 -14013 -33849 -13995
rect -33651 -14004 -33633 -13986
rect -31446 -13977 -31419 -13950
rect -31374 -13968 -31347 -13941
rect -31896 -14022 -31878 -14004
rect -31680 -14013 -31662 -13995
rect -33417 -14463 -33390 -14436
rect -33345 -14454 -33318 -14427
rect -31446 -14454 -31419 -14427
rect -31374 -14445 -31347 -14418
rect -33867 -14508 -33849 -14490
rect -33651 -14499 -33633 -14481
rect -31896 -14499 -31878 -14481
rect -31680 -14490 -31662 -14472
rect -31446 -14850 -31419 -14823
rect -31374 -14841 -31347 -14814
rect -31896 -14895 -31878 -14877
rect -31680 -14886 -31662 -14868
rect -33417 -14958 -33390 -14931
rect -33345 -14949 -33318 -14922
rect -33867 -15003 -33849 -14985
rect -33651 -14994 -33633 -14976
rect -31446 -15318 -31419 -15291
rect -31374 -15309 -31347 -15282
rect -33417 -15372 -33390 -15345
rect -33345 -15363 -33318 -15336
rect -31896 -15363 -31878 -15345
rect -31680 -15354 -31662 -15336
rect -33867 -15417 -33849 -15399
rect -33651 -15408 -33633 -15390
rect -33417 -15903 -33390 -15876
rect -33345 -15894 -33318 -15867
rect -33867 -15948 -33849 -15930
rect -33651 -15939 -33633 -15921
<< pdcontact >>
rect -30222 10296 -30186 10332
rect -30222 10224 -30186 10260
rect -30222 10125 -30186 10161
rect -29412 10296 -29376 10332
rect -30222 10053 -30186 10089
rect -30222 9936 -30186 9972
rect -30222 9855 -30186 9891
rect -30222 9774 -30186 9810
rect -30222 9693 -30186 9729
rect -29412 10224 -29376 10260
rect -29412 10125 -29376 10161
rect -28530 10296 -28494 10332
rect -29412 10053 -29376 10089
rect -29412 9936 -29376 9972
rect -29412 9855 -29376 9891
rect -29412 9774 -29376 9810
rect -29412 9693 -29376 9729
rect -28530 10224 -28494 10260
rect -28530 10125 -28494 10161
rect -28530 10053 -28494 10089
rect -28530 9936 -28494 9972
rect -28530 9855 -28494 9891
rect -28530 9774 -28494 9810
rect -28530 9693 -28494 9729
rect -30357 9315 -30339 9333
rect -30303 9306 -30285 9324
rect -30204 9315 -30186 9333
rect -30141 9315 -30123 9333
rect -29907 9351 -29880 9378
rect -29835 9342 -29808 9369
rect -29331 9378 -29313 9396
rect -29277 9369 -29259 9387
rect -29178 9378 -29160 9396
rect -29115 9378 -29097 9396
rect -28881 9414 -28854 9441
rect -28809 9405 -28782 9432
rect -29691 8955 -29673 8973
rect -29538 8946 -29520 8964
rect -29466 8955 -29448 8973
rect -29412 8946 -29394 8964
rect -30222 8199 -30186 8235
rect -30222 8127 -30186 8163
rect -30222 8028 -30186 8064
rect -29412 8199 -29376 8235
rect -30222 7956 -30186 7992
rect -30222 7839 -30186 7875
rect -30222 7758 -30186 7794
rect -30222 7677 -30186 7713
rect -30222 7596 -30186 7632
rect -29412 8127 -29376 8163
rect -29412 8028 -29376 8064
rect -28530 8199 -28494 8235
rect -29412 7956 -29376 7992
rect -29412 7839 -29376 7875
rect -29412 7758 -29376 7794
rect -29412 7677 -29376 7713
rect -29412 7596 -29376 7632
rect -28530 8127 -28494 8163
rect -28530 8028 -28494 8064
rect -28530 7956 -28494 7992
rect -28530 7839 -28494 7875
rect -28530 7758 -28494 7794
rect -28530 7677 -28494 7713
rect -28530 7596 -28494 7632
rect -30357 7218 -30339 7236
rect -30303 7209 -30285 7227
rect -30204 7218 -30186 7236
rect -30141 7218 -30123 7236
rect -29907 7254 -29880 7281
rect -29835 7245 -29808 7272
rect -29331 7281 -29313 7299
rect -29277 7272 -29259 7290
rect -29178 7281 -29160 7299
rect -29115 7281 -29097 7299
rect -28881 7317 -28854 7344
rect -28809 7308 -28782 7335
rect -29691 6858 -29673 6876
rect -29538 6849 -29520 6867
rect -29466 6858 -29448 6876
rect -29412 6849 -29394 6867
rect -30222 6084 -30186 6120
rect -30222 6012 -30186 6048
rect -30222 5913 -30186 5949
rect -29412 6084 -29376 6120
rect -30222 5841 -30186 5877
rect -30222 5724 -30186 5760
rect -30222 5643 -30186 5679
rect -30222 5562 -30186 5598
rect -30222 5481 -30186 5517
rect -29412 6012 -29376 6048
rect -29412 5913 -29376 5949
rect -28530 6084 -28494 6120
rect -29412 5841 -29376 5877
rect -29412 5724 -29376 5760
rect -29412 5643 -29376 5679
rect -29412 5562 -29376 5598
rect -29412 5481 -29376 5517
rect -28530 6012 -28494 6048
rect -28530 5913 -28494 5949
rect -28530 5841 -28494 5877
rect -28530 5724 -28494 5760
rect -28530 5643 -28494 5679
rect -28530 5562 -28494 5598
rect -28530 5481 -28494 5517
rect -30357 5103 -30339 5121
rect -30303 5094 -30285 5112
rect -30204 5103 -30186 5121
rect -30141 5103 -30123 5121
rect -29907 5139 -29880 5166
rect -29835 5130 -29808 5157
rect -29331 5166 -29313 5184
rect -29277 5157 -29259 5175
rect -29178 5166 -29160 5184
rect -29115 5166 -29097 5184
rect -28881 5202 -28854 5229
rect -28809 5193 -28782 5220
rect -29691 4743 -29673 4761
rect -29538 4734 -29520 4752
rect -29466 4743 -29448 4761
rect -29412 4734 -29394 4752
rect -30222 4149 -30186 4185
rect -30222 4077 -30186 4113
rect -30222 3978 -30186 4014
rect -29412 4149 -29376 4185
rect -30222 3906 -30186 3942
rect -30222 3789 -30186 3825
rect -30222 3708 -30186 3744
rect -30222 3627 -30186 3663
rect -30222 3546 -30186 3582
rect -29412 4077 -29376 4113
rect -29412 3978 -29376 4014
rect -28530 4149 -28494 4185
rect -29412 3906 -29376 3942
rect -29412 3789 -29376 3825
rect -29412 3708 -29376 3744
rect -29412 3627 -29376 3663
rect -29412 3546 -29376 3582
rect -28530 4077 -28494 4113
rect -28530 3978 -28494 4014
rect -28530 3906 -28494 3942
rect -28530 3789 -28494 3825
rect -28530 3708 -28494 3744
rect -28530 3627 -28494 3663
rect -28530 3546 -28494 3582
rect -30357 3168 -30339 3186
rect -30303 3159 -30285 3177
rect -30204 3168 -30186 3186
rect -30141 3168 -30123 3186
rect -29907 3204 -29880 3231
rect -29835 3195 -29808 3222
rect -29331 3231 -29313 3249
rect -29277 3222 -29259 3240
rect -29178 3231 -29160 3249
rect -29115 3231 -29097 3249
rect -28881 3267 -28854 3294
rect -28809 3258 -28782 3285
rect -29691 2808 -29673 2826
rect -29538 2799 -29520 2817
rect -29466 2808 -29448 2826
rect -29412 2799 -29394 2817
rect -29862 459 -29826 495
rect -29862 387 -29826 423
rect -29862 288 -29826 324
rect -29511 369 -29484 396
rect -29439 360 -29412 387
rect -29862 216 -29826 252
rect -29862 99 -29826 135
rect -29862 18 -29826 54
rect -29862 -63 -29826 -27
rect -29862 -144 -29826 -108
rect -28305 99 -28278 126
rect -29142 63 -29115 90
rect -29070 54 -29043 81
rect -28755 63 -28737 81
rect -28701 54 -28683 72
rect -28602 63 -28584 81
rect -28539 63 -28521 81
rect -28233 90 -28206 117
rect -33435 -315 -33408 -288
rect -33885 -351 -33867 -333
rect -33831 -360 -33813 -342
rect -33732 -351 -33714 -333
rect -33669 -351 -33651 -333
rect -33363 -324 -33336 -297
rect -29862 -486 -29826 -450
rect -33435 -810 -33408 -783
rect -33885 -846 -33867 -828
rect -33831 -855 -33813 -837
rect -33732 -846 -33714 -828
rect -33669 -846 -33651 -828
rect -33363 -819 -33336 -792
rect -34461 -1098 -34443 -1080
rect -34308 -1107 -34290 -1089
rect -34236 -1098 -34218 -1080
rect -34182 -1107 -34164 -1089
rect -33435 -1224 -33408 -1197
rect -33885 -1260 -33867 -1242
rect -33831 -1269 -33813 -1251
rect -33732 -1260 -33714 -1242
rect -33669 -1260 -33651 -1242
rect -33363 -1233 -33336 -1206
rect -33435 -1755 -33408 -1728
rect -33885 -1791 -33867 -1773
rect -33831 -1800 -33813 -1782
rect -33732 -1791 -33714 -1773
rect -33669 -1791 -33651 -1773
rect -33363 -1764 -33336 -1737
rect -33435 -2322 -33408 -2295
rect -33885 -2358 -33867 -2340
rect -33831 -2367 -33813 -2349
rect -33732 -2358 -33714 -2340
rect -33669 -2358 -33651 -2340
rect -33363 -2331 -33336 -2304
rect -33435 -2817 -33408 -2790
rect -33885 -2853 -33867 -2835
rect -33831 -2862 -33813 -2844
rect -33732 -2853 -33714 -2835
rect -33669 -2853 -33651 -2835
rect -33363 -2826 -33336 -2799
rect -33435 -3231 -33408 -3204
rect -33885 -3267 -33867 -3249
rect -33831 -3276 -33813 -3258
rect -33732 -3267 -33714 -3249
rect -33669 -3267 -33651 -3249
rect -33363 -3240 -33336 -3213
rect -33435 -3762 -33408 -3735
rect -33885 -3798 -33867 -3780
rect -33831 -3807 -33813 -3789
rect -33732 -3798 -33714 -3780
rect -33669 -3798 -33651 -3780
rect -33363 -3771 -33336 -3744
rect -33417 -8172 -33390 -8145
rect -33867 -8208 -33849 -8190
rect -33813 -8217 -33795 -8199
rect -33714 -8208 -33696 -8190
rect -33651 -8208 -33633 -8190
rect -33345 -8181 -33318 -8154
rect -29862 -558 -29826 -522
rect -29862 -657 -29826 -621
rect -29511 -576 -29484 -549
rect -29439 -585 -29412 -558
rect -29862 -729 -29826 -693
rect -28377 -711 -28350 -684
rect -29862 -846 -29826 -810
rect -29862 -927 -29826 -891
rect -29160 -747 -29133 -720
rect -29088 -756 -29061 -729
rect -28827 -747 -28809 -729
rect -28773 -756 -28755 -738
rect -28674 -747 -28656 -729
rect -28611 -747 -28593 -729
rect -28305 -720 -28278 -693
rect -27999 -747 -27981 -729
rect -27945 -756 -27927 -738
rect -27549 -711 -27522 -684
rect -27846 -747 -27828 -729
rect -27783 -747 -27765 -729
rect -27477 -720 -27450 -693
rect -27126 -756 -27108 -738
rect -26793 -765 -26775 -747
rect -26721 -756 -26703 -738
rect -26667 -765 -26649 -747
rect -29862 -1008 -29826 -972
rect -29862 -1089 -29826 -1053
rect -29862 -1503 -29826 -1467
rect -29862 -1575 -29826 -1539
rect -29862 -1674 -29826 -1638
rect -28674 -1530 -28647 -1503
rect -28611 -1539 -28584 -1512
rect -28548 -1530 -28521 -1503
rect -28485 -1539 -28458 -1512
rect -28404 -1530 -28377 -1503
rect -28341 -1539 -28314 -1512
rect -28278 -1530 -28251 -1503
rect -28215 -1539 -28188 -1512
rect -28152 -1530 -28125 -1503
rect -28080 -1539 -28053 -1512
rect -27882 -1521 -27855 -1494
rect -27819 -1539 -27792 -1512
rect -29511 -1593 -29484 -1566
rect -29439 -1602 -29412 -1575
rect -29178 -1593 -29151 -1566
rect -29106 -1602 -29079 -1575
rect -29862 -1746 -29826 -1710
rect -29862 -1863 -29826 -1827
rect -29862 -1944 -29826 -1908
rect -29862 -2025 -29826 -1989
rect -29862 -2106 -29826 -2070
rect -29862 -2799 -29826 -2763
rect -29862 -2871 -29826 -2835
rect -29862 -2970 -29826 -2934
rect -28827 -2826 -28800 -2799
rect -28764 -2835 -28737 -2808
rect -28701 -2826 -28674 -2799
rect -28638 -2835 -28611 -2808
rect -28557 -2826 -28530 -2799
rect -28494 -2835 -28467 -2808
rect -28431 -2826 -28404 -2799
rect -28368 -2835 -28341 -2808
rect -28305 -2826 -28278 -2799
rect -28233 -2835 -28206 -2808
rect -28035 -2817 -28008 -2790
rect -27972 -2835 -27945 -2808
rect -29511 -2889 -29484 -2862
rect -29439 -2898 -29412 -2871
rect -29232 -2889 -29205 -2862
rect -29160 -2898 -29133 -2871
rect -29862 -3042 -29826 -3006
rect -29862 -3159 -29826 -3123
rect -29862 -3240 -29826 -3204
rect -29862 -3321 -29826 -3285
rect -29862 -3402 -29826 -3366
rect -29862 -3870 -29826 -3834
rect -29862 -3942 -29826 -3906
rect -29862 -4041 -29826 -4005
rect -29511 -3960 -29484 -3933
rect -29439 -3969 -29412 -3942
rect -29862 -4113 -29826 -4077
rect -29862 -4230 -29826 -4194
rect -29862 -4311 -29826 -4275
rect -29862 -4392 -29826 -4356
rect -29862 -4473 -29826 -4437
rect -28305 -4230 -28278 -4203
rect -29142 -4266 -29115 -4239
rect -29070 -4275 -29043 -4248
rect -28755 -4266 -28737 -4248
rect -28701 -4275 -28683 -4257
rect -28602 -4266 -28584 -4248
rect -28539 -4266 -28521 -4248
rect -28233 -4239 -28206 -4212
rect -29862 -4815 -29826 -4779
rect -29862 -4887 -29826 -4851
rect -29862 -4986 -29826 -4950
rect -29511 -4905 -29484 -4878
rect -29439 -4914 -29412 -4887
rect -29862 -5058 -29826 -5022
rect -28377 -5040 -28350 -5013
rect -29862 -5175 -29826 -5139
rect -29862 -5256 -29826 -5220
rect -29160 -5076 -29133 -5049
rect -29088 -5085 -29061 -5058
rect -28827 -5076 -28809 -5058
rect -28773 -5085 -28755 -5067
rect -28674 -5076 -28656 -5058
rect -28611 -5076 -28593 -5058
rect -28305 -5049 -28278 -5022
rect -27999 -5076 -27981 -5058
rect -27945 -5085 -27927 -5067
rect -27549 -5040 -27522 -5013
rect -27846 -5076 -27828 -5058
rect -27783 -5076 -27765 -5058
rect -27477 -5049 -27450 -5022
rect -27126 -5085 -27108 -5067
rect -26793 -5094 -26775 -5076
rect -26721 -5085 -26703 -5067
rect -26667 -5094 -26649 -5076
rect -29862 -5337 -29826 -5301
rect -29862 -5418 -29826 -5382
rect -29862 -5832 -29826 -5796
rect -29862 -5904 -29826 -5868
rect -29862 -6003 -29826 -5967
rect -28674 -5859 -28647 -5832
rect -28611 -5868 -28584 -5841
rect -28548 -5859 -28521 -5832
rect -28485 -5868 -28458 -5841
rect -28404 -5859 -28377 -5832
rect -28341 -5868 -28314 -5841
rect -28278 -5859 -28251 -5832
rect -28215 -5868 -28188 -5841
rect -28152 -5859 -28125 -5832
rect -28080 -5868 -28053 -5841
rect -27882 -5850 -27855 -5823
rect -27819 -5868 -27792 -5841
rect -29511 -5922 -29484 -5895
rect -29439 -5931 -29412 -5904
rect -29178 -5922 -29151 -5895
rect -29106 -5931 -29079 -5904
rect -29862 -6075 -29826 -6039
rect -29862 -6192 -29826 -6156
rect -29862 -6273 -29826 -6237
rect -29862 -6354 -29826 -6318
rect -29862 -6435 -29826 -6399
rect -33417 -8667 -33390 -8640
rect -33867 -8703 -33849 -8685
rect -33813 -8712 -33795 -8694
rect -33714 -8703 -33696 -8685
rect -33651 -8703 -33633 -8685
rect -33345 -8676 -33318 -8649
rect -33417 -9081 -33390 -9054
rect -33867 -9117 -33849 -9099
rect -33813 -9126 -33795 -9108
rect -33714 -9117 -33696 -9099
rect -33651 -9117 -33633 -9099
rect -33345 -9090 -33318 -9063
rect -33417 -9612 -33390 -9585
rect -33867 -9648 -33849 -9630
rect -33813 -9657 -33795 -9639
rect -33714 -9648 -33696 -9630
rect -33651 -9648 -33633 -9630
rect -33345 -9621 -33318 -9594
rect -33417 -10089 -33390 -10062
rect -33867 -10125 -33849 -10107
rect -33813 -10134 -33795 -10116
rect -33714 -10125 -33696 -10107
rect -33651 -10125 -33633 -10107
rect -33345 -10098 -33318 -10071
rect -33417 -10584 -33390 -10557
rect -33867 -10620 -33849 -10602
rect -33813 -10629 -33795 -10611
rect -33714 -10620 -33696 -10602
rect -33651 -10620 -33633 -10602
rect -33345 -10593 -33318 -10566
rect -35415 -11511 -35388 -11484
rect -35865 -11547 -35847 -11529
rect -35811 -11556 -35793 -11538
rect -35712 -11547 -35694 -11529
rect -35649 -11547 -35631 -11529
rect -35343 -11520 -35316 -11493
rect -35415 -11979 -35388 -11952
rect -35865 -12015 -35847 -11997
rect -35811 -12024 -35793 -12006
rect -35712 -12015 -35694 -11997
rect -35649 -12015 -35631 -11997
rect -35343 -11988 -35316 -11961
rect -33417 -10998 -33390 -10971
rect -33867 -11034 -33849 -11016
rect -33813 -11043 -33795 -11025
rect -33714 -11034 -33696 -11016
rect -33651 -11034 -33633 -11016
rect -33345 -11007 -33318 -10980
rect -29862 -7128 -29826 -7092
rect -29862 -7200 -29826 -7164
rect -29862 -7299 -29826 -7263
rect -29511 -7218 -29484 -7191
rect -29439 -7227 -29412 -7200
rect -29862 -7371 -29826 -7335
rect -29862 -7488 -29826 -7452
rect -29862 -7569 -29826 -7533
rect -29862 -7650 -29826 -7614
rect -29862 -7731 -29826 -7695
rect -29862 -8667 -29826 -8631
rect -29862 -8739 -29826 -8703
rect -29862 -8838 -29826 -8802
rect -28827 -7155 -28800 -7128
rect -28764 -7164 -28737 -7137
rect -28701 -7155 -28674 -7128
rect -28638 -7164 -28611 -7137
rect -28557 -7155 -28530 -7128
rect -28494 -7164 -28467 -7137
rect -28431 -7155 -28404 -7128
rect -28368 -7164 -28341 -7137
rect -28305 -7155 -28278 -7128
rect -28233 -7164 -28206 -7137
rect -28035 -7146 -28008 -7119
rect -27972 -7164 -27945 -7137
rect -29232 -7218 -29205 -7191
rect -29160 -7227 -29133 -7200
rect -29511 -8757 -29484 -8730
rect -29439 -8766 -29412 -8739
rect -29862 -8910 -29826 -8874
rect -29862 -9027 -29826 -8991
rect -29862 -9108 -29826 -9072
rect -29862 -9189 -29826 -9153
rect -29862 -9270 -29826 -9234
rect -29862 -9612 -29826 -9576
rect -29862 -9684 -29826 -9648
rect -29862 -9783 -29826 -9747
rect -29511 -9702 -29484 -9675
rect -29439 -9711 -29412 -9684
rect -29862 -9855 -29826 -9819
rect -29862 -9972 -29826 -9936
rect -29862 -10053 -29826 -10017
rect -29862 -10134 -29826 -10098
rect -26406 -9765 -26379 -9738
rect -28206 -9810 -28179 -9783
rect -28143 -9819 -28116 -9792
rect -28080 -9810 -28053 -9783
rect -28017 -9819 -27990 -9792
rect -27936 -9810 -27909 -9783
rect -27873 -9819 -27846 -9792
rect -27810 -9810 -27783 -9783
rect -27747 -9819 -27720 -9792
rect -27684 -9810 -27657 -9783
rect -27612 -9819 -27585 -9792
rect -27414 -9801 -27387 -9774
rect -27351 -9819 -27324 -9792
rect -26856 -9801 -26838 -9783
rect -26802 -9810 -26784 -9792
rect -26703 -9801 -26685 -9783
rect -26640 -9801 -26622 -9783
rect -26334 -9774 -26307 -9747
rect -29862 -10215 -29826 -10179
rect -29862 -10629 -29826 -10593
rect -29862 -10701 -29826 -10665
rect -29862 -10800 -29826 -10764
rect -29511 -10719 -29484 -10692
rect -29439 -10728 -29412 -10701
rect -29862 -10872 -29826 -10836
rect -29862 -10989 -29826 -10953
rect -29862 -11070 -29826 -11034
rect -29862 -11151 -29826 -11115
rect -29862 -11232 -29826 -11196
rect -33417 -11529 -33390 -11502
rect -33867 -11565 -33849 -11547
rect -33813 -11574 -33795 -11556
rect -33714 -11565 -33696 -11547
rect -33651 -11565 -33633 -11547
rect -33345 -11538 -33318 -11511
rect -36207 -12168 -36180 -12141
rect -36135 -12177 -36108 -12150
rect -35415 -12420 -35388 -12393
rect -35865 -12456 -35847 -12438
rect -36198 -12492 -36171 -12465
rect -35811 -12465 -35793 -12447
rect -35712 -12456 -35694 -12438
rect -35649 -12456 -35631 -12438
rect -35343 -12429 -35316 -12402
rect -29862 -11925 -29826 -11889
rect -33417 -12393 -33390 -12366
rect -33867 -12429 -33849 -12411
rect -36126 -12501 -36099 -12474
rect -33813 -12438 -33795 -12420
rect -33714 -12429 -33696 -12411
rect -33651 -12429 -33633 -12411
rect -33345 -12402 -33318 -12375
rect -35415 -12834 -35388 -12807
rect -35865 -12870 -35847 -12852
rect -35811 -12879 -35793 -12861
rect -35712 -12870 -35694 -12852
rect -35649 -12870 -35631 -12852
rect -35343 -12843 -35316 -12816
rect -29862 -11997 -29826 -11961
rect -29862 -12096 -29826 -12060
rect -29511 -12015 -29484 -11988
rect -29439 -12024 -29412 -11997
rect -29862 -12168 -29826 -12132
rect -29862 -12285 -29826 -12249
rect -29862 -12366 -29826 -12330
rect -29862 -12447 -29826 -12411
rect -29862 -12528 -29826 -12492
rect -33417 -12888 -33390 -12861
rect -33867 -12924 -33849 -12906
rect -33813 -12933 -33795 -12915
rect -33714 -12924 -33696 -12906
rect -33651 -12924 -33633 -12906
rect -33345 -12897 -33318 -12870
rect -33417 -13302 -33390 -13275
rect -33867 -13338 -33849 -13320
rect -33813 -13347 -33795 -13329
rect -33714 -13338 -33696 -13320
rect -33651 -13338 -33633 -13320
rect -33345 -13311 -33318 -13284
rect -33417 -13833 -33390 -13806
rect -33867 -13869 -33849 -13851
rect -33813 -13878 -33795 -13860
rect -33714 -13869 -33696 -13851
rect -33651 -13869 -33633 -13851
rect -33345 -13842 -33318 -13815
rect -31446 -13842 -31419 -13815
rect -31896 -13878 -31878 -13860
rect -31842 -13887 -31824 -13869
rect -31743 -13878 -31725 -13860
rect -31680 -13878 -31662 -13860
rect -31374 -13851 -31347 -13824
rect -33417 -14328 -33390 -14301
rect -33867 -14364 -33849 -14346
rect -33813 -14373 -33795 -14355
rect -33714 -14364 -33696 -14346
rect -33651 -14364 -33633 -14346
rect -33345 -14337 -33318 -14310
rect -31446 -14319 -31419 -14292
rect -31896 -14355 -31878 -14337
rect -31842 -14364 -31824 -14346
rect -31743 -14355 -31725 -14337
rect -31680 -14355 -31662 -14337
rect -31374 -14328 -31347 -14301
rect -31446 -14715 -31419 -14688
rect -31896 -14751 -31878 -14733
rect -31842 -14760 -31824 -14742
rect -31743 -14751 -31725 -14733
rect -31680 -14751 -31662 -14733
rect -31374 -14724 -31347 -14697
rect -33417 -14823 -33390 -14796
rect -33867 -14859 -33849 -14841
rect -33813 -14868 -33795 -14850
rect -33714 -14859 -33696 -14841
rect -33651 -14859 -33633 -14841
rect -33345 -14832 -33318 -14805
rect -31446 -15183 -31419 -15156
rect -33417 -15237 -33390 -15210
rect -33867 -15273 -33849 -15255
rect -33813 -15282 -33795 -15264
rect -33714 -15273 -33696 -15255
rect -33651 -15273 -33633 -15255
rect -33345 -15246 -33318 -15219
rect -31896 -15219 -31878 -15201
rect -31842 -15228 -31824 -15210
rect -31743 -15219 -31725 -15201
rect -31680 -15219 -31662 -15201
rect -31374 -15192 -31347 -15165
rect -33417 -15768 -33390 -15741
rect -33867 -15804 -33849 -15786
rect -33813 -15813 -33795 -15795
rect -33714 -15804 -33696 -15786
rect -33651 -15804 -33633 -15786
rect -33345 -15777 -33318 -15750
<< psubstratepcontact >>
rect -30600 9900 -30564 9936
rect -30600 9810 -30564 9846
rect -29790 9900 -29754 9936
rect -29790 9810 -29754 9846
rect -28908 9900 -28872 9936
rect -28908 9810 -28872 9846
rect -30600 7803 -30564 7839
rect -30600 7713 -30564 7749
rect -29790 7803 -29754 7839
rect -29790 7713 -29754 7749
rect -28908 7803 -28872 7839
rect -28908 7713 -28872 7749
rect -30600 5688 -30564 5724
rect -30600 5598 -30564 5634
rect -29790 5688 -29754 5724
rect -29790 5598 -29754 5634
rect -28908 5688 -28872 5724
rect -28908 5598 -28872 5634
rect -30600 3753 -30564 3789
rect -30600 3663 -30564 3699
rect -29790 3753 -29754 3789
rect -29790 3663 -29754 3699
rect -28908 3753 -28872 3789
rect -28908 3663 -28872 3699
rect -30240 63 -30204 99
rect -30240 -27 -30204 9
rect -30240 -882 -30204 -846
rect -30240 -972 -30204 -936
rect -30240 -1899 -30204 -1863
rect -30240 -1989 -30204 -1953
rect -30240 -3195 -30204 -3159
rect -30240 -3285 -30204 -3249
rect -30240 -4266 -30204 -4230
rect -30240 -4356 -30204 -4320
rect -30240 -5211 -30204 -5175
rect -30240 -5301 -30204 -5265
rect -30240 -6228 -30204 -6192
rect -30240 -6318 -30204 -6282
rect -30240 -7524 -30204 -7488
rect -30240 -7614 -30204 -7578
rect -30240 -9063 -30204 -9027
rect -30240 -9153 -30204 -9117
rect -30240 -10008 -30204 -9972
rect -30240 -10098 -30204 -10062
rect -30240 -11025 -30204 -10989
rect -30240 -11115 -30204 -11079
rect -30240 -12321 -30204 -12285
rect -30240 -12411 -30204 -12375
<< nsubstratencontact >>
rect -30105 9900 -30069 9936
rect -30105 9810 -30069 9846
rect -29295 9900 -29259 9936
rect -29295 9810 -29259 9846
rect -28413 9900 -28377 9936
rect -28413 9810 -28377 9846
rect -30105 7803 -30069 7839
rect -30105 7713 -30069 7749
rect -29295 7803 -29259 7839
rect -29295 7713 -29259 7749
rect -28413 7803 -28377 7839
rect -28413 7713 -28377 7749
rect -30105 5688 -30069 5724
rect -30105 5598 -30069 5634
rect -29295 5688 -29259 5724
rect -29295 5598 -29259 5634
rect -28413 5688 -28377 5724
rect -28413 5598 -28377 5634
rect -30105 3753 -30069 3789
rect -30105 3663 -30069 3699
rect -29295 3753 -29259 3789
rect -29295 3663 -29259 3699
rect -28413 3753 -28377 3789
rect -28413 3663 -28377 3699
rect -29745 63 -29709 99
rect -29745 -27 -29709 9
rect -29745 -882 -29709 -846
rect -29745 -972 -29709 -936
rect -29745 -1899 -29709 -1863
rect -29745 -1989 -29709 -1953
rect -29745 -3195 -29709 -3159
rect -29745 -3285 -29709 -3249
rect -29745 -4266 -29709 -4230
rect -29745 -4356 -29709 -4320
rect -29745 -5211 -29709 -5175
rect -29745 -5301 -29709 -5265
rect -29745 -6228 -29709 -6192
rect -29745 -6318 -29709 -6282
rect -29745 -7524 -29709 -7488
rect -29745 -7614 -29709 -7578
rect -29745 -9063 -29709 -9027
rect -29745 -9153 -29709 -9117
rect -29745 -10008 -29709 -9972
rect -29745 -10098 -29709 -10062
rect -29745 -11025 -29709 -10989
rect -29745 -11115 -29709 -11079
rect -29745 -12321 -29709 -12285
rect -29745 -12411 -29709 -12375
<< polysilicon >>
rect -30537 10377 -30096 10395
rect -30537 10287 -30519 10377
rect -30690 10269 -30483 10287
rect -30429 10269 -30420 10287
rect -30402 10269 -30231 10287
rect -30168 10269 -30141 10287
rect -30852 7803 -30834 9882
rect -30690 9630 -30672 10269
rect -30402 10116 -30384 10269
rect -30114 10116 -30096 10377
rect -29727 10377 -29286 10395
rect -29727 10287 -29709 10377
rect -29880 10269 -29673 10287
rect -29619 10269 -29610 10287
rect -29592 10269 -29421 10287
rect -29358 10269 -29331 10287
rect -30051 10170 -29952 10188
rect -30645 10098 -30483 10116
rect -30429 10098 -30384 10116
rect -30267 10098 -30231 10116
rect -30168 10098 -30096 10116
rect -30645 9756 -30627 10098
rect -30357 9918 -30321 9945
rect -30546 9900 -30483 9918
rect -30429 9900 -30231 9918
rect -30168 9900 -30123 9918
rect -29970 9909 -29952 10170
rect -30348 9837 -30330 9900
rect -30024 9891 -29952 9909
rect -30519 9828 -30330 9837
rect -30357 9765 -30348 9801
rect -30330 9765 -30321 9801
rect -30357 9756 -30321 9765
rect -30645 9738 -30483 9756
rect -30429 9738 -30231 9756
rect -30168 9738 -30123 9756
rect -30690 9612 -30321 9630
rect -30024 9612 -30006 9891
rect -29970 9882 -29952 9891
rect -29952 9864 -29943 9882
rect -29880 9630 -29862 10269
rect -29592 10116 -29574 10269
rect -29304 10116 -29286 10377
rect -28845 10377 -28404 10395
rect -28845 10287 -28827 10377
rect -28998 10269 -28791 10287
rect -28737 10269 -28728 10287
rect -28710 10269 -28539 10287
rect -28476 10269 -28449 10287
rect -29241 10170 -29115 10188
rect -29835 10098 -29673 10116
rect -29619 10098 -29574 10116
rect -29457 10098 -29421 10116
rect -29358 10098 -29286 10116
rect -29835 9756 -29817 10098
rect -29547 9918 -29511 9945
rect -29736 9900 -29673 9918
rect -29619 9900 -29421 9918
rect -29358 9900 -29313 9918
rect -29538 9837 -29520 9900
rect -29133 9882 -29115 10170
rect -29133 9864 -29088 9882
rect -29691 9828 -29520 9837
rect -29547 9765 -29511 9801
rect -29547 9756 -29538 9765
rect -29835 9738 -29673 9756
rect -29619 9738 -29538 9756
rect -29520 9756 -29511 9765
rect -29520 9738 -29421 9756
rect -29358 9738 -29313 9756
rect -29880 9612 -29511 9630
rect -30159 9594 -30006 9612
rect -30159 9486 -30141 9594
rect -29484 9531 -29466 9738
rect -29133 9549 -29115 9864
rect -29070 9864 -29052 9882
rect -28998 9630 -28980 10269
rect -28710 10116 -28692 10269
rect -28422 10116 -28404 10377
rect -28359 10161 -28278 10197
rect -28953 10098 -28791 10116
rect -28737 10098 -28692 10116
rect -28575 10098 -28539 10116
rect -28476 10098 -28404 10116
rect -28953 9756 -28935 10098
rect -28665 9918 -28629 9945
rect -28854 9900 -28791 9918
rect -28737 9900 -28539 9918
rect -28476 9900 -28431 9918
rect -28656 9837 -28638 9900
rect -28809 9828 -28638 9837
rect -28665 9792 -28629 9801
rect -28665 9765 -28656 9792
rect -28638 9765 -28629 9792
rect -28665 9756 -28629 9765
rect -28953 9738 -28791 9756
rect -28737 9738 -28539 9756
rect -28476 9738 -28431 9756
rect -28998 9612 -28629 9630
rect -28602 9594 -28584 9738
rect -28494 9639 -28179 9657
rect -30429 9468 -30141 9486
rect -30051 9513 -29466 9531
rect -29403 9531 -29115 9549
rect -29025 9576 -28584 9594
rect -30429 9234 -30411 9468
rect -30330 9342 -30312 9369
rect -30168 9342 -30150 9369
rect -30330 9234 -30312 9297
rect -30429 9216 -30312 9234
rect -30330 9198 -30312 9216
rect -30168 9225 -30150 9297
rect -30051 9225 -30033 9513
rect -29871 9378 -29853 9495
rect -29871 9288 -29853 9324
rect -29862 9261 -29853 9288
rect -29871 9252 -29853 9261
rect -30168 9207 -30033 9225
rect -29871 9207 -29853 9225
rect -30168 9198 -30150 9207
rect -30330 9162 -30312 9171
rect -30168 9162 -30150 9171
rect -29772 8892 -29754 9297
rect -29610 9027 -29592 9432
rect -29529 9189 -29511 9477
rect -29403 9297 -29385 9531
rect -29304 9405 -29286 9432
rect -29142 9405 -29124 9432
rect -29304 9297 -29286 9360
rect -29403 9279 -29286 9297
rect -29304 9261 -29286 9279
rect -29142 9288 -29124 9360
rect -29025 9288 -29007 9576
rect -29142 9270 -29007 9288
rect -29142 9261 -29124 9270
rect -29304 9225 -29286 9234
rect -29142 9225 -29124 9234
rect -28989 9216 -28971 9549
rect -28845 9441 -28827 9558
rect -28845 9351 -28827 9387
rect -28836 9324 -28827 9351
rect -28746 9333 -28710 9360
rect -28845 9315 -28827 9324
rect -28845 9270 -28827 9288
rect -28728 9144 -28710 9333
rect -29502 9126 -28710 9144
rect -29655 8982 -29637 9000
rect -29565 8982 -29547 9000
rect -29655 8892 -29637 8937
rect -29772 8874 -29637 8892
rect -29655 8847 -29637 8874
rect -29565 8865 -29547 8937
rect -29502 8865 -29484 9126
rect -29439 8982 -29421 9000
rect -29565 8856 -29484 8865
rect -29439 8892 -29421 8937
rect -29430 8874 -29421 8892
rect -29565 8847 -29547 8856
rect -29439 8847 -29421 8874
rect -29655 8811 -29637 8820
rect -29565 8811 -29547 8820
rect -29439 8811 -29421 8820
rect -28197 8343 -28179 9639
rect -28197 8316 -27765 8343
rect -30537 8280 -30096 8298
rect -30537 8190 -30519 8280
rect -30852 6507 -30834 7785
rect -30690 8172 -30483 8190
rect -30429 8172 -30420 8190
rect -30402 8172 -30231 8190
rect -30168 8172 -30141 8190
rect -30690 7533 -30672 8172
rect -30402 8019 -30384 8172
rect -30114 8019 -30096 8280
rect -29727 8280 -29286 8298
rect -29727 8190 -29709 8280
rect -29880 8172 -29673 8190
rect -29619 8172 -29610 8190
rect -29592 8172 -29421 8190
rect -29358 8172 -29331 8190
rect -30051 8073 -29952 8091
rect -30645 8001 -30483 8019
rect -30429 8001 -30384 8019
rect -30267 8001 -30231 8019
rect -30168 8001 -30096 8019
rect -30645 7659 -30627 8001
rect -30357 7821 -30321 7848
rect -30546 7803 -30483 7821
rect -30429 7803 -30231 7821
rect -30168 7803 -30123 7821
rect -29970 7812 -29952 8073
rect -30348 7740 -30330 7803
rect -30024 7794 -29952 7812
rect -30528 7731 -30330 7740
rect -30357 7677 -30348 7704
rect -30330 7677 -30321 7704
rect -30357 7659 -30321 7677
rect -30645 7641 -30483 7659
rect -30429 7641 -30231 7659
rect -30168 7641 -30123 7659
rect -30690 7515 -30321 7533
rect -30024 7515 -30006 7794
rect -29970 7785 -29952 7794
rect -29952 7767 -29943 7785
rect -29880 7533 -29862 8172
rect -29592 8019 -29574 8172
rect -29304 8019 -29286 8280
rect -28845 8280 -28404 8298
rect -28845 8190 -28827 8280
rect -28998 8172 -28791 8190
rect -28737 8172 -28728 8190
rect -28710 8172 -28539 8190
rect -28476 8172 -28449 8190
rect -29241 8073 -29115 8091
rect -29835 8001 -29673 8019
rect -29619 8001 -29574 8019
rect -29457 8001 -29421 8019
rect -29358 8001 -29286 8019
rect -29835 7659 -29817 8001
rect -29547 7821 -29511 7848
rect -29736 7803 -29673 7821
rect -29619 7803 -29421 7821
rect -29358 7803 -29313 7821
rect -29538 7740 -29520 7803
rect -29133 7785 -29115 8073
rect -29133 7767 -29088 7785
rect -29691 7731 -29520 7740
rect -29547 7668 -29511 7704
rect -29547 7659 -29538 7668
rect -29835 7641 -29673 7659
rect -29619 7641 -29538 7659
rect -29520 7659 -29511 7668
rect -29520 7641 -29421 7659
rect -29358 7641 -29313 7659
rect -29880 7515 -29511 7533
rect -30159 7497 -30006 7515
rect -30159 7389 -30141 7497
rect -29484 7434 -29466 7641
rect -29133 7452 -29115 7767
rect -29070 7767 -29052 7785
rect -28998 7533 -28980 8172
rect -28710 8019 -28692 8172
rect -28422 8019 -28404 8280
rect -28359 8064 -28278 8100
rect -28953 8001 -28791 8019
rect -28737 8001 -28692 8019
rect -28575 8001 -28539 8019
rect -28476 8001 -28404 8019
rect -28953 7659 -28935 8001
rect -28665 7821 -28629 7848
rect -28854 7803 -28791 7821
rect -28737 7803 -28539 7821
rect -28476 7803 -28431 7821
rect -28656 7740 -28638 7803
rect -28809 7731 -28638 7740
rect -28665 7677 -28656 7704
rect -28638 7677 -28629 7704
rect -28665 7659 -28629 7677
rect -28953 7641 -28791 7659
rect -28737 7641 -28539 7659
rect -28476 7641 -28431 7659
rect -28998 7515 -28629 7533
rect -28602 7497 -28584 7641
rect -28485 7551 -27909 7569
rect -30429 7371 -30141 7389
rect -30051 7416 -29466 7434
rect -29403 7434 -29115 7452
rect -29025 7479 -28584 7497
rect -30429 7137 -30411 7371
rect -30330 7245 -30312 7272
rect -30168 7245 -30150 7272
rect -30330 7137 -30312 7200
rect -30429 7119 -30312 7137
rect -30330 7101 -30312 7119
rect -30168 7128 -30150 7200
rect -30051 7128 -30033 7416
rect -29871 7281 -29853 7398
rect -29871 7191 -29853 7227
rect -29862 7164 -29853 7191
rect -29871 7155 -29853 7164
rect -30168 7110 -30033 7128
rect -29871 7110 -29853 7128
rect -30168 7101 -30150 7110
rect -30330 7065 -30312 7074
rect -30168 7065 -30150 7074
rect -29772 6795 -29754 7200
rect -29610 6930 -29592 7335
rect -29529 7092 -29511 7380
rect -29403 7200 -29385 7434
rect -29304 7308 -29286 7335
rect -29142 7308 -29124 7335
rect -29304 7200 -29286 7263
rect -29403 7182 -29286 7200
rect -29304 7164 -29286 7182
rect -29142 7191 -29124 7263
rect -29025 7191 -29007 7479
rect -29142 7173 -29007 7191
rect -29142 7164 -29124 7173
rect -29304 7128 -29286 7137
rect -29142 7128 -29124 7137
rect -28989 7119 -28971 7452
rect -28845 7344 -28827 7461
rect -28845 7254 -28827 7290
rect -28836 7227 -28827 7254
rect -28746 7236 -28710 7263
rect -28845 7218 -28827 7227
rect -28845 7173 -28827 7191
rect -28728 7047 -28710 7236
rect -29502 7029 -28710 7047
rect -29655 6885 -29637 6903
rect -29565 6885 -29547 6903
rect -29655 6795 -29637 6840
rect -29772 6777 -29637 6795
rect -29655 6750 -29637 6777
rect -29565 6768 -29547 6840
rect -29502 6768 -29484 7029
rect -29439 6885 -29421 6903
rect -29565 6759 -29484 6768
rect -29439 6795 -29421 6840
rect -29430 6777 -29421 6795
rect -29565 6750 -29547 6759
rect -29439 6750 -29421 6777
rect -29655 6714 -29637 6723
rect -29565 6714 -29547 6723
rect -29439 6714 -29421 6723
rect -36801 6480 -30834 6507
rect -36801 1152 -36783 6480
rect -30852 5688 -30834 6480
rect -30537 6165 -30096 6183
rect -30537 6075 -30519 6165
rect -30852 4833 -30834 5670
rect -30690 6057 -30483 6075
rect -30429 6057 -30420 6075
rect -30402 6057 -30231 6075
rect -30168 6057 -30141 6075
rect -30690 5418 -30672 6057
rect -30402 5904 -30384 6057
rect -30114 5904 -30096 6165
rect -29727 6165 -29286 6183
rect -29727 6075 -29709 6165
rect -29880 6057 -29673 6075
rect -29619 6057 -29610 6075
rect -29592 6057 -29421 6075
rect -29358 6057 -29331 6075
rect -30051 5958 -29952 5976
rect -30645 5886 -30483 5904
rect -30429 5886 -30384 5904
rect -30267 5886 -30231 5904
rect -30168 5886 -30096 5904
rect -30645 5544 -30627 5886
rect -30357 5706 -30321 5733
rect -30546 5688 -30483 5706
rect -30429 5688 -30231 5706
rect -30168 5688 -30123 5706
rect -29970 5697 -29952 5958
rect -30348 5625 -30330 5688
rect -30024 5679 -29952 5697
rect -30528 5616 -30330 5625
rect -30357 5553 -30348 5589
rect -30330 5553 -30321 5589
rect -30357 5544 -30321 5553
rect -30645 5526 -30483 5544
rect -30429 5526 -30231 5544
rect -30168 5526 -30123 5544
rect -30690 5400 -30321 5418
rect -30024 5400 -30006 5679
rect -29970 5670 -29952 5679
rect -29952 5652 -29943 5670
rect -29880 5418 -29862 6057
rect -29592 5904 -29574 6057
rect -29304 5904 -29286 6165
rect -28845 6165 -28404 6183
rect -28845 6075 -28827 6165
rect -28998 6057 -28791 6075
rect -28737 6057 -28728 6075
rect -28710 6057 -28539 6075
rect -28476 6057 -28449 6075
rect -29241 5958 -29115 5976
rect -29835 5886 -29673 5904
rect -29619 5886 -29574 5904
rect -29457 5886 -29421 5904
rect -29358 5886 -29286 5904
rect -29835 5544 -29817 5886
rect -29547 5706 -29511 5733
rect -29736 5688 -29673 5706
rect -29619 5688 -29421 5706
rect -29358 5688 -29313 5706
rect -29538 5625 -29520 5688
rect -29133 5670 -29115 5958
rect -29133 5652 -29088 5670
rect -29691 5616 -29520 5625
rect -29547 5553 -29511 5589
rect -29547 5544 -29538 5553
rect -29835 5526 -29673 5544
rect -29619 5526 -29538 5544
rect -29511 5526 -29421 5544
rect -29358 5526 -29313 5544
rect -29880 5400 -29511 5418
rect -30159 5382 -30006 5400
rect -30159 5274 -30141 5382
rect -29484 5319 -29466 5526
rect -29133 5337 -29115 5652
rect -29070 5652 -29052 5670
rect -28998 5418 -28980 6057
rect -28710 5904 -28692 6057
rect -28422 5904 -28404 6165
rect -28359 5949 -28278 5985
rect -28953 5886 -28791 5904
rect -28737 5886 -28692 5904
rect -28575 5886 -28539 5904
rect -28476 5886 -28404 5904
rect -28953 5544 -28935 5886
rect -28665 5706 -28629 5733
rect -28854 5688 -28791 5706
rect -28737 5688 -28539 5706
rect -28476 5688 -28431 5706
rect -28656 5625 -28638 5688
rect -28809 5616 -28638 5625
rect -28665 5580 -28629 5589
rect -28665 5562 -28656 5580
rect -28638 5562 -28629 5580
rect -28665 5544 -28629 5562
rect -28953 5526 -28791 5544
rect -28737 5526 -28539 5544
rect -28476 5526 -28431 5544
rect -28998 5400 -28629 5418
rect -28602 5382 -28584 5526
rect -30429 5256 -30141 5274
rect -30051 5301 -29466 5319
rect -29403 5319 -29115 5337
rect -29025 5364 -28584 5382
rect -30429 5022 -30411 5256
rect -30330 5130 -30312 5157
rect -30168 5130 -30150 5157
rect -30330 5022 -30312 5085
rect -30429 5004 -30312 5022
rect -30330 4986 -30312 5004
rect -30168 5013 -30150 5085
rect -30051 5013 -30033 5301
rect -29871 5166 -29853 5283
rect -29871 5076 -29853 5112
rect -29862 5049 -29853 5076
rect -29871 5040 -29853 5049
rect -30168 4995 -30033 5013
rect -29871 4995 -29853 5013
rect -30168 4986 -30150 4995
rect -30330 4950 -30312 4959
rect -30168 4950 -30150 4959
rect -30852 4815 -30708 4833
rect -30726 3825 -30708 4815
rect -29772 4680 -29754 5085
rect -29610 4815 -29592 5220
rect -29529 4977 -29511 5265
rect -29403 5085 -29385 5319
rect -29304 5193 -29286 5220
rect -29142 5193 -29124 5220
rect -29304 5085 -29286 5148
rect -29403 5067 -29286 5085
rect -29304 5049 -29286 5067
rect -29142 5076 -29124 5148
rect -29025 5076 -29007 5364
rect -29142 5058 -29007 5076
rect -29142 5049 -29124 5058
rect -29304 5013 -29286 5022
rect -29142 5013 -29124 5022
rect -28989 5004 -28971 5337
rect -28845 5229 -28827 5346
rect -28845 5139 -28827 5175
rect -28836 5112 -28827 5139
rect -28746 5121 -28710 5148
rect -28845 5103 -28827 5112
rect -28845 5058 -28827 5076
rect -28728 4932 -28710 5121
rect -29502 4914 -28710 4932
rect -29655 4770 -29637 4788
rect -29565 4770 -29547 4788
rect -29655 4680 -29637 4725
rect -29772 4662 -29637 4680
rect -29655 4635 -29637 4662
rect -29565 4653 -29547 4725
rect -29502 4653 -29484 4914
rect -29439 4770 -29421 4788
rect -29565 4644 -29484 4653
rect -29439 4680 -29421 4725
rect -27927 4680 -27909 7551
rect -27783 6795 -27765 8316
rect -29430 4662 -29421 4680
rect -29367 4662 -27909 4680
rect -29565 4635 -29547 4644
rect -29439 4635 -29421 4662
rect -29655 4599 -29637 4608
rect -29565 4599 -29547 4608
rect -29439 4599 -29421 4608
rect -30537 4230 -30096 4248
rect -30537 4140 -30519 4230
rect -30726 3789 -30708 3807
rect -30690 4122 -30483 4140
rect -30429 4122 -30420 4140
rect -30402 4122 -30231 4140
rect -30168 4122 -30141 4140
rect -30690 3483 -30672 4122
rect -30402 3969 -30384 4122
rect -30114 3969 -30096 4230
rect -29727 4230 -29286 4248
rect -29727 4140 -29709 4230
rect -29880 4122 -29673 4140
rect -29619 4122 -29610 4140
rect -29592 4122 -29421 4140
rect -29358 4122 -29331 4140
rect -30051 4023 -29952 4041
rect -30645 3951 -30483 3969
rect -30429 3951 -30384 3969
rect -30267 3951 -30231 3969
rect -30168 3951 -30096 3969
rect -30645 3609 -30627 3951
rect -30357 3771 -30321 3798
rect -30546 3753 -30483 3771
rect -30429 3753 -30231 3771
rect -30168 3753 -30123 3771
rect -29970 3762 -29952 4023
rect -30528 3690 -30510 3726
rect -30348 3690 -30330 3753
rect -30024 3744 -29952 3762
rect -30528 3681 -30330 3690
rect -30357 3627 -30348 3654
rect -30330 3627 -30321 3654
rect -30357 3609 -30321 3627
rect -30645 3591 -30483 3609
rect -30429 3591 -30231 3609
rect -30168 3591 -30123 3609
rect -30690 3465 -30321 3483
rect -30024 3465 -30006 3744
rect -29970 3735 -29952 3744
rect -29952 3717 -29943 3735
rect -29880 3483 -29862 4122
rect -29592 3969 -29574 4122
rect -29304 3969 -29286 4230
rect -28845 4230 -28404 4248
rect -28845 4140 -28827 4230
rect -28998 4122 -28791 4140
rect -28737 4122 -28728 4140
rect -28710 4122 -28539 4140
rect -28476 4122 -28449 4140
rect -29241 4023 -29115 4041
rect -29835 3951 -29673 3969
rect -29619 3951 -29574 3969
rect -29457 3951 -29421 3969
rect -29358 3951 -29286 3969
rect -29835 3609 -29817 3951
rect -29547 3771 -29511 3798
rect -29736 3753 -29673 3771
rect -29619 3753 -29421 3771
rect -29358 3753 -29313 3771
rect -29538 3690 -29520 3753
rect -29133 3735 -29115 4023
rect -29133 3717 -29088 3735
rect -29691 3681 -29520 3690
rect -29547 3618 -29511 3654
rect -29547 3609 -29538 3618
rect -29835 3591 -29673 3609
rect -29619 3591 -29538 3609
rect -29511 3591 -29421 3609
rect -29358 3591 -29313 3609
rect -29880 3465 -29511 3483
rect -30159 3447 -30006 3465
rect -30159 3339 -30141 3447
rect -29484 3384 -29466 3591
rect -29133 3402 -29115 3717
rect -29070 3717 -29052 3735
rect -28998 3483 -28980 4122
rect -28710 3969 -28692 4122
rect -28422 3969 -28404 4230
rect -28359 4014 -28278 4050
rect -28953 3951 -28791 3969
rect -28737 3951 -28692 3969
rect -28575 3951 -28539 3969
rect -28476 3951 -28404 3969
rect -28953 3609 -28935 3951
rect -28665 3771 -28629 3798
rect -28854 3753 -28791 3771
rect -28737 3753 -28539 3771
rect -28476 3753 -28431 3771
rect -28656 3690 -28638 3753
rect -28809 3681 -28638 3690
rect -28665 3645 -28629 3654
rect -28665 3627 -28656 3645
rect -28638 3627 -28629 3645
rect -28665 3609 -28629 3627
rect -28953 3591 -28791 3609
rect -28737 3591 -28539 3609
rect -28476 3591 -28431 3609
rect -28998 3465 -28629 3483
rect -28602 3447 -28584 3591
rect -30429 3321 -30141 3339
rect -30051 3366 -29466 3384
rect -29403 3384 -29115 3402
rect -29025 3429 -28584 3447
rect -30429 3087 -30411 3321
rect -30330 3195 -30312 3222
rect -30168 3195 -30150 3222
rect -30330 3087 -30312 3150
rect -30429 3069 -30312 3087
rect -30330 3051 -30312 3069
rect -30168 3078 -30150 3150
rect -30051 3078 -30033 3366
rect -29871 3231 -29853 3348
rect -29871 3141 -29853 3177
rect -29862 3114 -29853 3141
rect -29871 3105 -29853 3114
rect -30168 3060 -30033 3078
rect -29871 3060 -29853 3078
rect -30168 3051 -30150 3060
rect -30330 3015 -30312 3024
rect -30168 3015 -30150 3024
rect -29772 2745 -29754 3150
rect -29610 2880 -29592 3285
rect -29529 3042 -29511 3330
rect -29403 3150 -29385 3384
rect -29304 3258 -29286 3285
rect -29142 3258 -29124 3285
rect -29304 3150 -29286 3213
rect -29403 3132 -29286 3150
rect -29304 3114 -29286 3132
rect -29142 3141 -29124 3213
rect -29025 3141 -29007 3429
rect -29142 3123 -29007 3141
rect -29142 3114 -29124 3123
rect -29304 3078 -29286 3087
rect -29142 3078 -29124 3087
rect -28989 3069 -28971 3402
rect -28845 3294 -28827 3411
rect -28845 3204 -28827 3240
rect -28836 3177 -28827 3204
rect -28746 3186 -28710 3213
rect -28845 3168 -28827 3177
rect -28845 3123 -28827 3141
rect -28728 2997 -28710 3186
rect -29502 2979 -28710 2997
rect -29655 2835 -29637 2853
rect -29565 2835 -29547 2853
rect -29655 2745 -29637 2790
rect -29772 2727 -29637 2745
rect -29655 2700 -29637 2727
rect -29565 2718 -29547 2790
rect -29502 2718 -29484 2979
rect -29439 2835 -29421 2853
rect -29565 2709 -29484 2718
rect -29439 2745 -29421 2790
rect -29430 2727 -29421 2745
rect -29565 2700 -29547 2709
rect -29439 2700 -29421 2727
rect -29655 2664 -29637 2673
rect -29565 2664 -29547 2673
rect -29439 2664 -29421 2673
rect -30177 540 -29736 558
rect -28350 549 -28332 3348
rect -30177 450 -30159 540
rect -30330 432 -30123 450
rect -30069 432 -30060 450
rect -30042 432 -29871 450
rect -29808 432 -29781 450
rect -30699 -99 -30366 -81
rect -33399 -288 -33381 -171
rect -30330 -207 -30312 432
rect -30042 279 -30024 432
rect -29754 279 -29736 540
rect -28422 531 -28332 549
rect -29475 396 -29457 414
rect -29475 306 -29457 342
rect -30285 261 -30123 279
rect -30069 261 -30024 279
rect -29907 261 -29871 279
rect -29808 261 -29736 279
rect -29691 279 -29511 306
rect -29466 279 -29457 306
rect -29475 270 -29457 279
rect -30285 -81 -30267 261
rect -29475 225 -29457 243
rect -29997 81 -29961 108
rect -30177 63 -30168 81
rect -30141 63 -30123 81
rect -30069 63 -29871 81
rect -29808 63 -29763 81
rect -29988 -9 -29970 63
rect -29997 -81 -29961 -36
rect -30249 -99 -30123 -81
rect -30069 -99 -29871 -81
rect -29808 -99 -29763 -81
rect -30330 -225 -29961 -207
rect -29781 -288 -29763 -99
rect -29439 -99 -29421 189
rect -28422 153 -28404 531
rect -28269 126 -28251 243
rect -29106 90 -29088 108
rect -28728 90 -28710 117
rect -28566 90 -28548 117
rect -29106 0 -29088 36
rect -28728 9 -28710 45
rect -29097 -27 -29088 0
rect -29016 -18 -28710 9
rect -29106 -36 -29088 -27
rect -28728 -54 -28710 -18
rect -28566 -27 -28548 45
rect -28269 36 -28251 72
rect -28260 9 -28251 36
rect -28269 0 -28251 9
rect -28620 -45 -28548 -27
rect -28269 -45 -28251 -27
rect -28620 -54 -28611 -45
rect -28566 -54 -28548 -45
rect -29106 -81 -29088 -63
rect -28728 -90 -28710 -81
rect -29439 -117 -29151 -99
rect -28620 -288 -28611 -81
rect -28566 -90 -28548 -81
rect -33858 -324 -33840 -297
rect -33696 -324 -33678 -297
rect -29781 -306 -28611 -288
rect -33858 -432 -33840 -369
rect -34029 -450 -33840 -432
rect -34029 -927 -34011 -450
rect -33858 -468 -33840 -450
rect -33696 -468 -33678 -369
rect -33399 -378 -33381 -342
rect -33390 -405 -33381 -378
rect -33399 -414 -33381 -405
rect -30177 -405 -29736 -387
rect -33399 -459 -33381 -441
rect -30177 -495 -30159 -405
rect -33858 -504 -33840 -495
rect -33696 -549 -33678 -495
rect -30330 -513 -30123 -495
rect -30069 -513 -30060 -495
rect -30042 -513 -29871 -495
rect -29808 -513 -29781 -495
rect -33858 -819 -33840 -792
rect -33696 -819 -33678 -747
rect -33399 -783 -33381 -666
rect -33858 -927 -33840 -864
rect -34029 -945 -33840 -927
rect -34425 -1071 -34407 -1053
rect -34335 -1071 -34317 -1053
rect -34209 -1071 -34191 -1053
rect -34425 -1206 -34407 -1116
rect -34335 -1206 -34317 -1116
rect -34209 -1161 -34191 -1116
rect -34029 -1161 -34011 -945
rect -33858 -963 -33840 -945
rect -33696 -963 -33678 -864
rect -33399 -873 -33381 -837
rect -33390 -900 -33381 -873
rect -33399 -909 -33381 -900
rect -33399 -954 -33381 -936
rect -33858 -999 -33840 -990
rect -33696 -999 -33678 -990
rect -30879 -1044 -30366 -1026
rect -34200 -1179 -34191 -1161
rect -34119 -1179 -34011 -1161
rect -34209 -1206 -34191 -1179
rect -36918 -1278 -35820 -1269
rect -34425 -1278 -34407 -1233
rect -36918 -1305 -34407 -1278
rect -36918 -11052 -36900 -1305
rect -34335 -1341 -34317 -1233
rect -34209 -1242 -34191 -1233
rect -36783 -1377 -34317 -1341
rect -34029 -1350 -34011 -1179
rect -33399 -1197 -33381 -1080
rect -33858 -1233 -33840 -1206
rect -33696 -1233 -33678 -1206
rect -33858 -1350 -33840 -1278
rect -34029 -1368 -33840 -1350
rect -36801 -10737 -36783 -1413
rect -34029 -1872 -34011 -1368
rect -33858 -1377 -33840 -1368
rect -33696 -1377 -33678 -1278
rect -33399 -1287 -33381 -1251
rect -33390 -1314 -33381 -1287
rect -33399 -1323 -33381 -1314
rect -33399 -1368 -33381 -1350
rect -33858 -1413 -33840 -1404
rect -33696 -1458 -33678 -1404
rect -33399 -1728 -33381 -1611
rect -33858 -1764 -33840 -1737
rect -33696 -1764 -33678 -1737
rect -33858 -1872 -33840 -1809
rect -34029 -1890 -33840 -1872
rect -34029 -2439 -34011 -1890
rect -33858 -1908 -33840 -1890
rect -33696 -1908 -33678 -1809
rect -33399 -1818 -33381 -1782
rect -33390 -1845 -33381 -1818
rect -33399 -1854 -33381 -1845
rect -33399 -1899 -33381 -1881
rect -33858 -1944 -33840 -1935
rect -33696 -1989 -33678 -1935
rect -33399 -2295 -33381 -2178
rect -33858 -2331 -33840 -2304
rect -33696 -2331 -33678 -2304
rect -33858 -2439 -33840 -2376
rect -34029 -2457 -33840 -2439
rect -34029 -2934 -34011 -2457
rect -33858 -2475 -33840 -2457
rect -33696 -2475 -33678 -2376
rect -33399 -2385 -33381 -2349
rect -33390 -2412 -33381 -2385
rect -33399 -2421 -33381 -2412
rect -33399 -2466 -33381 -2448
rect -33858 -2511 -33840 -2502
rect -33696 -2547 -33678 -2502
rect -33399 -2790 -33381 -2673
rect -33858 -2826 -33840 -2799
rect -33696 -2826 -33678 -2799
rect -33858 -2934 -33840 -2871
rect -34029 -2952 -33840 -2934
rect -34029 -3357 -34011 -2952
rect -33858 -2970 -33840 -2952
rect -33696 -2970 -33678 -2871
rect -33399 -2880 -33381 -2844
rect -33390 -2907 -33381 -2880
rect -33399 -2916 -33381 -2907
rect -33399 -2961 -33381 -2943
rect -33858 -3006 -33840 -2997
rect -33696 -3051 -33678 -2997
rect -33399 -3204 -33381 -3087
rect -33858 -3240 -33840 -3213
rect -33696 -3240 -33678 -3213
rect -33858 -3357 -33840 -3285
rect -34029 -3375 -33840 -3357
rect -34029 -3879 -34011 -3375
rect -33858 -3384 -33840 -3375
rect -33696 -3384 -33678 -3285
rect -33399 -3294 -33381 -3258
rect -33390 -3321 -33381 -3294
rect -33399 -3330 -33381 -3321
rect -33399 -3375 -33381 -3357
rect -33858 -3420 -33840 -3411
rect -33696 -3474 -33678 -3411
rect -33399 -3735 -33381 -3618
rect -33858 -3771 -33840 -3744
rect -33696 -3771 -33678 -3744
rect -31167 -3744 -31023 -3726
rect -33858 -3879 -33840 -3816
rect -34029 -3897 -33840 -3879
rect -33858 -3915 -33840 -3897
rect -33696 -3915 -33678 -3816
rect -33399 -3825 -33381 -3789
rect -33390 -3852 -33381 -3825
rect -33399 -3861 -33381 -3852
rect -33399 -3906 -33381 -3888
rect -33858 -3951 -33840 -3942
rect -33696 -3987 -33678 -3942
rect -33381 -8145 -33363 -8028
rect -33840 -8181 -33822 -8154
rect -33678 -8181 -33660 -8154
rect -33840 -8289 -33822 -8226
rect -34011 -8307 -33822 -8289
rect -34011 -8784 -33993 -8307
rect -33840 -8325 -33822 -8307
rect -33678 -8325 -33660 -8226
rect -33381 -8235 -33363 -8199
rect -31284 -8226 -31266 -6723
rect -31167 -7902 -31149 -3744
rect -30960 -5373 -30942 -1053
rect -30330 -1152 -30312 -513
rect -30042 -666 -30024 -513
rect -29754 -666 -29736 -405
rect -29475 -549 -29457 -531
rect -29475 -639 -29457 -603
rect -30285 -684 -30123 -666
rect -30069 -684 -30024 -666
rect -29907 -684 -29871 -666
rect -29808 -684 -29736 -666
rect -29691 -666 -29511 -639
rect -29466 -666 -29457 -639
rect -29475 -675 -29457 -666
rect -30285 -1026 -30267 -684
rect -28341 -684 -28323 -567
rect -29475 -720 -29457 -702
rect -29124 -720 -29106 -702
rect -28800 -720 -28782 -693
rect -28638 -720 -28620 -693
rect -29997 -864 -29961 -837
rect -30132 -882 -30123 -864
rect -30069 -882 -29871 -864
rect -29808 -882 -29763 -864
rect -29988 -954 -29970 -882
rect -29475 -909 -29457 -756
rect -27972 -720 -27954 -693
rect -29124 -810 -29106 -774
rect -28800 -801 -28782 -765
rect -29115 -837 -29106 -810
rect -29016 -828 -28782 -801
rect -29124 -846 -29106 -837
rect -28800 -864 -28782 -828
rect -28638 -837 -28620 -765
rect -28341 -774 -28323 -738
rect -28332 -801 -28323 -774
rect -28242 -792 -28125 -765
rect -28341 -810 -28323 -801
rect -28152 -801 -28125 -792
rect -27972 -801 -27954 -765
rect -28692 -855 -28620 -837
rect -28152 -828 -27954 -801
rect -28341 -855 -28323 -837
rect -28692 -864 -28683 -855
rect -28638 -864 -28620 -855
rect -27972 -864 -27954 -828
rect -27882 -837 -27864 -576
rect -27513 -684 -27495 -567
rect -27810 -720 -27792 -693
rect -27090 -729 -27072 -711
rect -27036 -729 -27018 18
rect -27000 -729 -26982 -711
rect -26910 -729 -26892 -711
rect -26820 -729 -26802 -711
rect -26694 -729 -26676 -711
rect -27810 -837 -27792 -765
rect -27513 -774 -27495 -738
rect -27504 -801 -27495 -774
rect -27513 -810 -27495 -801
rect -27090 -801 -27072 -774
rect -27882 -855 -27792 -837
rect -27036 -801 -27018 -774
rect -27000 -801 -26982 -774
rect -26910 -792 -26892 -774
rect -27036 -819 -26982 -801
rect -27513 -855 -27495 -837
rect -27810 -864 -27792 -855
rect -27090 -864 -27072 -819
rect -27000 -864 -26982 -819
rect -26910 -864 -26892 -810
rect -26820 -792 -26802 -774
rect -26820 -864 -26802 -810
rect -26694 -819 -26676 -774
rect -26685 -837 -26676 -819
rect -26694 -864 -26676 -837
rect -29124 -891 -29106 -873
rect -28800 -900 -28782 -891
rect -29475 -927 -29169 -909
rect -29997 -1026 -29961 -981
rect -28692 -1026 -28683 -891
rect -28638 -900 -28620 -891
rect -27972 -900 -27954 -891
rect -27810 -900 -27792 -891
rect -27090 -900 -27072 -891
rect -27000 -900 -26982 -891
rect -26910 -900 -26892 -891
rect -26820 -900 -26802 -891
rect -26694 -900 -26676 -891
rect -30249 -1044 -30123 -1026
rect -30069 -1044 -29871 -1026
rect -29808 -1044 -28683 -1026
rect -30330 -1170 -29961 -1152
rect -30177 -1422 -29736 -1404
rect -30177 -1512 -30159 -1422
rect -30330 -1530 -30123 -1512
rect -30069 -1530 -30060 -1512
rect -30042 -1530 -29871 -1512
rect -29808 -1530 -29781 -1512
rect -30888 -2061 -30366 -2043
rect -30330 -2169 -30312 -1530
rect -30042 -1683 -30024 -1530
rect -29754 -1683 -29736 -1422
rect -28638 -1494 -28620 -1485
rect -28512 -1494 -28494 -1485
rect -28368 -1494 -28350 -1485
rect -28242 -1494 -28224 -1485
rect -28107 -1494 -28089 -1485
rect -27846 -1494 -27828 -1485
rect -29475 -1566 -29457 -1548
rect -29142 -1566 -29124 -1548
rect -28638 -1602 -28620 -1548
rect -29475 -1656 -29457 -1620
rect -29142 -1656 -29124 -1620
rect -28629 -1629 -28620 -1602
rect -28512 -1620 -28494 -1548
rect -28368 -1620 -28350 -1548
rect -28242 -1620 -28224 -1548
rect -28107 -1620 -28089 -1548
rect -27846 -1584 -27828 -1548
rect -30285 -1701 -30123 -1683
rect -30069 -1701 -30024 -1683
rect -29907 -1701 -29871 -1683
rect -29808 -1701 -29736 -1683
rect -29691 -1683 -29511 -1656
rect -29466 -1683 -29457 -1656
rect -29133 -1683 -29124 -1656
rect -28638 -1674 -28620 -1629
rect -28512 -1674 -28494 -1647
rect -28368 -1674 -28350 -1647
rect -28242 -1674 -28224 -1647
rect -28107 -1674 -28089 -1647
rect -27846 -1674 -27828 -1611
rect -29475 -1692 -29457 -1683
rect -29142 -1692 -29124 -1683
rect -30285 -2043 -30267 -1701
rect -29475 -1737 -29457 -1719
rect -28638 -1710 -28620 -1701
rect -28512 -1710 -28494 -1701
rect -28368 -1710 -28350 -1701
rect -28242 -1710 -28224 -1701
rect -28107 -1710 -28089 -1701
rect -27846 -1710 -27828 -1701
rect -29142 -1737 -29124 -1719
rect -29421 -1773 -29178 -1755
rect -29142 -1773 -29133 -1755
rect -29997 -1881 -29961 -1854
rect -30186 -1899 -30123 -1881
rect -30069 -1899 -29871 -1881
rect -29808 -1899 -29763 -1881
rect -29943 -1962 -29925 -1899
rect -29997 -2007 -29961 -1998
rect -29997 -2034 -29988 -2007
rect -29970 -2034 -29961 -2007
rect -29997 -2043 -29961 -2034
rect -30249 -2061 -30123 -2043
rect -30069 -2061 -29871 -2043
rect -29808 -2061 -29763 -2043
rect -30330 -2187 -29961 -2169
rect -29916 -2322 -29898 -2196
rect -30735 -2340 -29898 -2322
rect -30177 -2718 -29736 -2700
rect -30177 -2808 -30159 -2718
rect -30330 -2826 -30123 -2808
rect -30069 -2826 -30060 -2808
rect -30042 -2826 -29871 -2808
rect -29808 -2826 -29781 -2808
rect -30330 -3465 -30312 -2826
rect -30042 -2979 -30024 -2826
rect -29754 -2979 -29736 -2718
rect -28791 -2790 -28773 -2781
rect -28665 -2790 -28647 -2781
rect -28521 -2790 -28503 -2781
rect -28395 -2790 -28377 -2781
rect -28260 -2790 -28242 -2781
rect -27999 -2790 -27981 -2781
rect -29475 -2862 -29457 -2844
rect -29196 -2862 -29178 -2844
rect -28791 -2898 -28773 -2844
rect -29475 -2952 -29457 -2916
rect -29196 -2952 -29178 -2916
rect -28782 -2925 -28773 -2898
rect -28665 -2916 -28647 -2844
rect -28521 -2916 -28503 -2844
rect -28395 -2916 -28377 -2844
rect -28260 -2916 -28242 -2844
rect -27999 -2880 -27981 -2844
rect -30285 -2997 -30123 -2979
rect -30069 -2997 -30024 -2979
rect -29907 -2997 -29871 -2979
rect -29808 -2997 -29736 -2979
rect -29691 -2979 -29511 -2952
rect -29466 -2979 -29457 -2952
rect -29187 -2979 -29178 -2952
rect -28791 -2970 -28773 -2925
rect -28665 -2970 -28647 -2943
rect -28521 -2970 -28503 -2943
rect -28395 -2970 -28377 -2943
rect -28260 -2970 -28242 -2943
rect -27999 -2970 -27981 -2907
rect -29475 -2988 -29457 -2979
rect -29196 -2988 -29178 -2979
rect -30285 -3339 -30267 -2997
rect -29475 -3033 -29457 -3015
rect -28791 -3006 -28773 -2997
rect -28665 -3006 -28647 -2997
rect -28521 -3006 -28503 -2997
rect -28395 -3006 -28377 -2997
rect -28260 -3006 -28242 -2997
rect -27999 -3006 -27981 -2997
rect -29196 -3033 -29178 -3015
rect -29997 -3177 -29961 -3150
rect -30186 -3195 -30123 -3177
rect -30069 -3195 -29871 -3177
rect -29808 -3195 -29763 -3177
rect -29943 -3249 -29925 -3195
rect -29997 -3303 -29961 -3294
rect -29997 -3321 -29988 -3303
rect -29970 -3321 -29961 -3303
rect -29997 -3339 -29961 -3321
rect -30285 -3357 -30123 -3339
rect -30069 -3357 -29871 -3339
rect -29808 -3357 -29763 -3339
rect -30330 -3483 -29961 -3465
rect -30177 -3789 -29736 -3771
rect -30177 -3879 -30159 -3789
rect -30330 -3897 -30123 -3879
rect -30069 -3897 -30060 -3879
rect -30042 -3897 -29871 -3879
rect -29808 -3897 -29781 -3879
rect -30330 -4536 -30312 -3897
rect -30042 -4050 -30024 -3897
rect -29754 -4050 -29736 -3789
rect -29610 -3861 -29583 -3240
rect -29475 -3933 -29457 -3915
rect -29475 -4023 -29457 -3987
rect -30285 -4068 -30123 -4050
rect -30069 -4068 -30024 -4050
rect -29907 -4068 -29871 -4050
rect -29808 -4068 -29736 -4050
rect -29691 -4050 -29511 -4023
rect -29466 -4050 -29457 -4023
rect -29475 -4059 -29457 -4050
rect -30285 -4410 -30267 -4068
rect -29475 -4104 -29457 -4086
rect -29997 -4248 -29961 -4221
rect -30186 -4266 -30123 -4248
rect -30069 -4266 -29871 -4248
rect -29808 -4266 -29763 -4248
rect -29988 -4338 -29970 -4266
rect -29997 -4410 -29961 -4365
rect -30285 -4428 -30123 -4410
rect -30069 -4428 -29871 -4410
rect -29808 -4428 -29763 -4410
rect -30330 -4554 -29961 -4536
rect -29781 -4617 -29763 -4428
rect -29439 -4428 -29421 -4140
rect -28269 -4203 -28251 -4086
rect -29106 -4239 -29088 -4221
rect -28728 -4239 -28710 -4212
rect -28566 -4239 -28548 -4212
rect -29106 -4329 -29088 -4293
rect -28728 -4320 -28710 -4284
rect -29097 -4356 -29088 -4329
rect -29016 -4347 -28710 -4320
rect -29106 -4365 -29088 -4356
rect -28728 -4383 -28710 -4347
rect -28566 -4356 -28548 -4284
rect -28269 -4293 -28251 -4257
rect -28260 -4320 -28251 -4293
rect -28269 -4329 -28251 -4320
rect -28620 -4374 -28548 -4356
rect -28269 -4374 -28251 -4356
rect -28620 -4383 -28611 -4374
rect -28566 -4383 -28548 -4374
rect -29106 -4410 -29088 -4392
rect -28728 -4419 -28710 -4410
rect -29439 -4446 -29151 -4428
rect -28620 -4617 -28611 -4410
rect -28566 -4419 -28548 -4410
rect -29781 -4635 -28611 -4617
rect -29781 -4662 -29763 -4635
rect -30780 -4680 -29763 -4662
rect -30177 -4734 -29736 -4716
rect -30177 -4824 -30159 -4734
rect -30330 -4842 -30123 -4824
rect -30069 -4842 -30060 -4824
rect -30042 -4842 -29871 -4824
rect -29808 -4842 -29781 -4824
rect -30330 -5481 -30312 -4842
rect -30042 -4995 -30024 -4842
rect -29754 -4995 -29736 -4734
rect -29475 -4878 -29457 -4860
rect -29475 -4968 -29457 -4932
rect -30285 -5013 -30123 -4995
rect -30069 -5013 -30024 -4995
rect -29907 -5013 -29871 -4995
rect -29808 -5013 -29736 -4995
rect -29691 -4995 -29511 -4968
rect -29466 -4995 -29457 -4968
rect -29475 -5004 -29457 -4995
rect -30285 -5355 -30267 -5013
rect -28341 -5013 -28323 -4896
rect -29475 -5049 -29457 -5031
rect -29124 -5049 -29106 -5031
rect -28800 -5049 -28782 -5022
rect -28638 -5049 -28620 -5022
rect -29997 -5193 -29961 -5166
rect -30186 -5211 -30123 -5193
rect -30069 -5211 -29871 -5193
rect -29808 -5211 -29763 -5193
rect -29988 -5283 -29970 -5211
rect -29475 -5238 -29457 -5085
rect -27972 -5049 -27954 -5022
rect -29124 -5139 -29106 -5103
rect -28800 -5130 -28782 -5094
rect -29115 -5166 -29106 -5139
rect -29016 -5157 -28782 -5130
rect -29124 -5175 -29106 -5166
rect -28800 -5193 -28782 -5157
rect -28638 -5166 -28620 -5094
rect -28341 -5103 -28323 -5067
rect -28332 -5130 -28323 -5103
rect -28242 -5121 -28125 -5094
rect -28341 -5139 -28323 -5130
rect -28152 -5130 -28125 -5121
rect -27972 -5130 -27954 -5094
rect -28692 -5184 -28620 -5166
rect -28152 -5157 -27954 -5130
rect -28341 -5184 -28323 -5166
rect -28692 -5193 -28683 -5184
rect -28638 -5193 -28620 -5184
rect -27972 -5193 -27954 -5157
rect -27882 -5166 -27864 -4905
rect -27513 -5013 -27495 -4896
rect -27810 -5049 -27792 -5022
rect -27090 -5058 -27072 -5040
rect -27036 -5058 -27018 -4311
rect -27000 -5058 -26982 -5040
rect -26910 -5058 -26892 -5040
rect -26820 -5058 -26802 -5040
rect -26694 -5058 -26676 -5040
rect -27810 -5166 -27792 -5094
rect -27513 -5103 -27495 -5067
rect -27504 -5130 -27495 -5103
rect -27513 -5139 -27495 -5130
rect -27090 -5130 -27072 -5103
rect -27882 -5184 -27792 -5166
rect -27036 -5130 -27018 -5103
rect -27000 -5130 -26982 -5103
rect -26910 -5121 -26892 -5103
rect -27036 -5148 -26982 -5130
rect -27513 -5184 -27495 -5166
rect -27810 -5193 -27792 -5184
rect -27090 -5193 -27072 -5148
rect -27000 -5193 -26982 -5148
rect -26910 -5193 -26892 -5139
rect -26820 -5121 -26802 -5103
rect -26820 -5193 -26802 -5139
rect -26694 -5148 -26676 -5103
rect -26685 -5166 -26676 -5148
rect -26694 -5193 -26676 -5166
rect -29124 -5220 -29106 -5202
rect -28800 -5229 -28782 -5220
rect -29475 -5256 -29169 -5238
rect -29997 -5355 -29961 -5310
rect -28692 -5355 -28683 -5220
rect -28638 -5229 -28620 -5220
rect -27972 -5229 -27954 -5220
rect -27810 -5229 -27792 -5220
rect -27090 -5229 -27072 -5220
rect -27000 -5229 -26982 -5220
rect -26910 -5229 -26892 -5220
rect -26820 -5229 -26802 -5220
rect -26694 -5229 -26676 -5220
rect -30285 -5373 -30240 -5355
rect -30213 -5373 -30123 -5355
rect -30069 -5373 -29871 -5355
rect -29808 -5373 -28683 -5355
rect -30330 -5499 -29961 -5481
rect -30240 -5670 -30213 -5526
rect -31086 -5688 -30213 -5670
rect -30177 -5751 -29736 -5733
rect -30177 -5841 -30159 -5751
rect -30330 -5859 -30123 -5841
rect -30069 -5859 -30060 -5841
rect -30042 -5859 -29871 -5841
rect -29808 -5859 -29781 -5841
rect -30330 -6498 -30312 -5859
rect -30042 -6012 -30024 -5859
rect -29754 -6012 -29736 -5751
rect -28638 -5823 -28620 -5814
rect -28512 -5823 -28494 -5814
rect -28368 -5823 -28350 -5814
rect -28242 -5823 -28224 -5814
rect -28107 -5823 -28089 -5814
rect -27846 -5823 -27828 -5814
rect -29475 -5895 -29457 -5877
rect -29142 -5895 -29124 -5877
rect -28638 -5931 -28620 -5877
rect -29475 -5985 -29457 -5949
rect -29142 -5985 -29124 -5949
rect -28629 -5958 -28620 -5931
rect -28512 -5949 -28494 -5877
rect -28368 -5949 -28350 -5877
rect -28242 -5949 -28224 -5877
rect -28107 -5949 -28089 -5877
rect -27846 -5913 -27828 -5877
rect -30285 -6030 -30123 -6012
rect -30069 -6030 -30024 -6012
rect -29907 -6030 -29871 -6012
rect -29808 -6030 -29736 -6012
rect -29691 -6012 -29511 -5985
rect -29466 -6012 -29457 -5985
rect -29133 -6012 -29124 -5985
rect -28638 -6003 -28620 -5958
rect -28512 -6003 -28494 -5976
rect -28368 -6003 -28350 -5976
rect -28242 -6003 -28224 -5976
rect -28107 -6003 -28089 -5976
rect -27846 -6003 -27828 -5940
rect -29475 -6021 -29457 -6012
rect -29142 -6021 -29124 -6012
rect -30285 -6372 -30267 -6030
rect -29475 -6066 -29457 -6048
rect -28638 -6039 -28620 -6030
rect -28512 -6039 -28494 -6030
rect -28368 -6039 -28350 -6030
rect -28242 -6039 -28224 -6030
rect -28107 -6039 -28089 -6030
rect -27846 -6039 -27828 -6030
rect -29142 -6066 -29124 -6048
rect -29421 -6102 -29178 -6084
rect -29142 -6102 -29133 -6084
rect -29997 -6210 -29961 -6183
rect -30186 -6228 -30123 -6210
rect -30069 -6228 -29871 -6210
rect -29808 -6228 -29763 -6210
rect -29943 -6291 -29925 -6228
rect -29997 -6336 -29961 -6327
rect -29997 -6363 -29988 -6336
rect -29970 -6363 -29961 -6336
rect -29997 -6372 -29961 -6363
rect -30285 -6390 -30240 -6372
rect -30222 -6390 -30123 -6372
rect -30069 -6390 -29871 -6372
rect -29808 -6390 -29763 -6372
rect -30330 -6516 -29961 -6498
rect -31077 -6651 -31050 -6642
rect -29943 -6651 -29925 -6534
rect -31077 -6669 -29925 -6651
rect -33372 -8262 -33363 -8235
rect -33291 -8253 -31266 -8226
rect -33336 -8262 -31266 -8253
rect -33381 -8271 -33363 -8262
rect -33381 -8316 -33363 -8298
rect -33840 -8361 -33822 -8352
rect -33678 -8406 -33660 -8352
rect -33381 -8640 -33363 -8523
rect -33840 -8676 -33822 -8649
rect -33678 -8676 -33660 -8649
rect -33840 -8784 -33822 -8721
rect -34011 -8802 -33822 -8784
rect -34011 -9207 -33993 -8802
rect -33840 -8820 -33822 -8802
rect -33678 -8820 -33660 -8721
rect -33381 -8730 -33363 -8694
rect -33372 -8757 -33363 -8730
rect -33291 -8748 -31545 -8721
rect -33381 -8766 -33363 -8757
rect -33381 -8811 -33363 -8793
rect -33840 -8856 -33822 -8847
rect -33678 -8901 -33660 -8847
rect -33381 -9054 -33363 -8937
rect -33840 -9090 -33822 -9063
rect -33678 -9090 -33660 -9063
rect -33840 -9207 -33822 -9135
rect -34011 -9225 -33822 -9207
rect -34011 -9729 -33993 -9225
rect -33840 -9234 -33822 -9225
rect -33678 -9234 -33660 -9135
rect -33381 -9144 -33363 -9108
rect -33372 -9171 -33363 -9144
rect -33291 -9153 -31437 -9135
rect -33381 -9180 -33363 -9171
rect -33381 -9225 -33363 -9207
rect -33840 -9270 -33822 -9261
rect -33678 -9315 -33660 -9261
rect -31284 -9387 -31266 -8262
rect -33381 -9585 -33363 -9468
rect -33840 -9621 -33822 -9594
rect -33678 -9621 -33660 -9594
rect -33840 -9729 -33822 -9666
rect -34011 -9747 -33822 -9729
rect -34011 -10206 -33993 -9747
rect -33840 -9765 -33822 -9747
rect -33678 -9765 -33660 -9666
rect -33381 -9675 -33363 -9639
rect -33372 -9702 -33363 -9675
rect -33291 -9693 -31437 -9666
rect -33381 -9711 -33363 -9702
rect -33381 -9756 -33363 -9738
rect -33840 -9801 -33822 -9792
rect -33678 -9855 -33660 -9792
rect -33381 -10062 -33363 -9945
rect -33840 -10098 -33822 -10071
rect -33678 -10098 -33660 -10071
rect -33840 -10206 -33822 -10143
rect -34011 -10224 -33822 -10206
rect -34011 -10701 -33993 -10224
rect -33840 -10242 -33822 -10224
rect -33678 -10242 -33660 -10143
rect -33381 -10152 -33363 -10116
rect -33372 -10179 -33363 -10152
rect -33291 -10170 -31491 -10143
rect -33381 -10188 -33363 -10179
rect -33381 -10233 -33363 -10215
rect -33840 -10278 -33822 -10269
rect -33678 -10332 -33660 -10269
rect -33381 -10557 -33363 -10440
rect -31518 -10449 -31491 -10170
rect -31518 -10467 -31455 -10449
rect -33840 -10593 -33822 -10566
rect -33678 -10593 -33660 -10566
rect -33840 -10701 -33822 -10638
rect -34011 -10719 -33822 -10701
rect -36801 -10773 -34866 -10737
rect -36918 -11070 -35082 -11052
rect -35379 -11484 -35361 -11367
rect -35838 -11520 -35820 -11493
rect -35676 -11520 -35658 -11493
rect -35838 -11619 -35820 -11565
rect -35676 -11637 -35658 -11565
rect -35379 -11574 -35361 -11538
rect -35100 -11565 -35082 -11070
rect -35370 -11601 -35361 -11574
rect -35289 -11592 -35082 -11565
rect -35379 -11610 -35361 -11601
rect -35838 -11664 -35820 -11637
rect -35379 -11655 -35361 -11637
rect -35676 -11664 -35658 -11655
rect -35838 -11700 -35820 -11691
rect -35676 -11700 -35658 -11691
rect -36306 -11952 -35910 -11934
rect -35379 -11952 -35361 -11835
rect -36306 -12231 -36288 -11952
rect -35928 -12096 -35910 -11952
rect -35838 -11988 -35820 -11961
rect -35676 -11988 -35658 -11961
rect -35838 -12096 -35820 -12033
rect -35928 -12114 -35820 -12096
rect -36171 -12141 -36153 -12123
rect -35838 -12132 -35820 -12114
rect -35676 -12105 -35658 -12033
rect -35379 -12042 -35361 -12006
rect -34884 -12033 -34866 -10773
rect -35370 -12069 -35361 -12042
rect -35289 -12060 -34866 -12033
rect -34011 -11124 -33993 -10719
rect -33840 -10737 -33822 -10719
rect -33678 -10737 -33660 -10638
rect -33381 -10647 -33363 -10611
rect -33372 -10674 -33363 -10647
rect -33291 -10665 -31518 -10638
rect -33381 -10683 -33363 -10674
rect -33381 -10728 -33363 -10710
rect -33840 -10773 -33822 -10764
rect -33678 -10818 -33660 -10764
rect -33381 -10971 -33363 -10854
rect -33840 -11007 -33822 -10980
rect -33678 -11007 -33660 -10980
rect -33840 -11124 -33822 -11052
rect -34011 -11142 -33822 -11124
rect -34011 -11646 -33993 -11142
rect -33840 -11151 -33822 -11142
rect -33678 -11151 -33660 -11052
rect -33381 -11061 -33363 -11025
rect -31077 -11052 -31050 -6669
rect -30960 -10602 -30942 -10368
rect -33372 -11088 -33363 -11061
rect -33291 -11079 -31050 -11052
rect -33381 -11097 -33363 -11088
rect -33381 -11142 -33363 -11124
rect -33840 -11187 -33822 -11178
rect -33678 -11232 -33660 -11178
rect -33381 -11502 -33363 -11385
rect -31077 -11403 -31050 -11079
rect -30879 -11169 -30861 -7065
rect -30177 -7047 -29736 -7029
rect -30177 -7137 -30159 -7047
rect -30330 -7155 -30123 -7137
rect -30069 -7155 -30060 -7137
rect -30042 -7155 -29871 -7137
rect -29808 -7155 -29781 -7137
rect -30330 -7794 -30312 -7155
rect -30042 -7308 -30024 -7155
rect -29754 -7308 -29736 -7047
rect -28791 -7119 -28773 -7110
rect -28665 -7119 -28647 -7110
rect -28521 -7119 -28503 -7110
rect -28395 -7119 -28377 -7110
rect -28260 -7119 -28242 -7110
rect -27999 -7119 -27981 -7110
rect -29475 -7191 -29457 -7173
rect -29475 -7281 -29457 -7245
rect -30285 -7326 -30123 -7308
rect -30069 -7326 -30024 -7308
rect -29907 -7326 -29871 -7308
rect -29808 -7326 -29736 -7308
rect -29691 -7308 -29511 -7281
rect -29466 -7308 -29457 -7281
rect -29475 -7317 -29457 -7308
rect -30285 -7668 -30267 -7326
rect -29475 -7362 -29457 -7344
rect -29997 -7506 -29961 -7479
rect -30186 -7524 -30123 -7506
rect -30069 -7524 -29871 -7506
rect -29808 -7524 -29763 -7506
rect -29943 -7578 -29925 -7524
rect -29997 -7632 -29961 -7623
rect -29997 -7650 -29988 -7632
rect -29970 -7650 -29961 -7632
rect -29997 -7668 -29961 -7650
rect -30285 -7686 -30123 -7668
rect -30069 -7686 -29871 -7668
rect -29808 -7686 -29763 -7668
rect -30330 -7812 -29961 -7794
rect -30177 -8586 -29736 -8568
rect -30177 -8676 -30159 -8586
rect -30330 -8694 -30123 -8676
rect -30069 -8694 -30060 -8676
rect -30042 -8694 -29871 -8676
rect -29808 -8694 -29781 -8676
rect -30330 -9333 -30312 -8694
rect -30042 -8847 -30024 -8694
rect -29754 -8847 -29736 -8586
rect -29340 -8631 -29322 -7137
rect -29196 -7191 -29178 -7173
rect -28791 -7227 -28773 -7173
rect -29196 -7281 -29178 -7245
rect -28782 -7254 -28773 -7227
rect -28665 -7245 -28647 -7173
rect -28521 -7245 -28503 -7173
rect -28395 -7245 -28377 -7173
rect -28260 -7245 -28242 -7173
rect -27999 -7209 -27981 -7173
rect -29187 -7308 -29178 -7281
rect -28791 -7299 -28773 -7254
rect -28665 -7299 -28647 -7272
rect -28521 -7299 -28503 -7272
rect -28395 -7299 -28377 -7272
rect -28260 -7299 -28242 -7272
rect -27999 -7299 -27981 -7236
rect -29196 -7317 -29178 -7308
rect -28791 -7335 -28773 -7326
rect -28665 -7335 -28647 -7326
rect -28521 -7335 -28503 -7326
rect -28395 -7335 -28377 -7326
rect -28260 -7335 -28242 -7326
rect -27999 -7335 -27981 -7326
rect -29196 -7362 -29178 -7344
rect -29475 -8730 -29457 -8712
rect -29475 -8820 -29457 -8784
rect -30285 -8865 -30123 -8847
rect -30069 -8865 -30024 -8847
rect -29907 -8865 -29871 -8847
rect -29808 -8865 -29736 -8847
rect -29691 -8847 -29511 -8820
rect -29466 -8847 -29457 -8820
rect -29385 -8838 -28899 -8811
rect -29475 -8856 -29457 -8847
rect -30285 -9207 -30267 -8865
rect -29475 -8901 -29457 -8883
rect -29997 -9045 -29961 -9018
rect -30168 -9063 -30123 -9045
rect -30069 -9063 -29871 -9045
rect -29808 -9063 -29763 -9045
rect -29997 -9207 -29961 -9162
rect -30285 -9225 -30123 -9207
rect -30069 -9225 -29871 -9207
rect -29808 -9225 -29763 -9207
rect -30330 -9351 -29961 -9333
rect -29781 -9432 -29763 -9225
rect -30177 -9531 -29736 -9513
rect -30177 -9621 -30159 -9531
rect -30330 -9639 -30123 -9621
rect -30069 -9639 -30060 -9621
rect -30042 -9639 -29871 -9621
rect -29808 -9639 -29781 -9621
rect -30330 -10278 -30312 -9639
rect -30042 -9792 -30024 -9639
rect -29754 -9792 -29736 -9531
rect -29475 -9675 -29457 -9657
rect -29475 -9765 -29457 -9729
rect -30285 -9810 -30123 -9792
rect -30069 -9810 -30024 -9792
rect -29907 -9810 -29871 -9792
rect -29808 -9810 -29736 -9792
rect -29691 -9792 -29511 -9765
rect -29466 -9792 -29457 -9765
rect -29385 -9783 -28998 -9756
rect -29475 -9801 -29457 -9792
rect -30285 -10152 -30267 -9810
rect -29475 -9846 -29457 -9828
rect -29997 -9990 -29961 -9963
rect -30168 -10008 -30123 -9990
rect -30069 -10008 -29871 -9990
rect -29808 -10008 -29763 -9990
rect -29997 -10152 -29961 -10107
rect -29016 -10107 -28998 -9783
rect -28926 -9882 -28899 -8838
rect -26370 -9738 -26352 -9621
rect -28170 -9774 -28152 -9765
rect -28044 -9774 -28026 -9765
rect -27900 -9774 -27882 -9765
rect -27774 -9774 -27756 -9765
rect -27639 -9774 -27621 -9765
rect -27378 -9774 -27360 -9765
rect -26829 -9774 -26811 -9747
rect -26667 -9774 -26649 -9747
rect -28170 -9882 -28152 -9828
rect -28926 -9909 -28152 -9882
rect -28170 -9954 -28152 -9909
rect -28044 -9954 -28026 -9828
rect -27900 -9954 -27882 -9828
rect -27774 -9954 -27756 -9828
rect -27639 -9954 -27621 -9828
rect -27378 -9864 -27360 -9828
rect -26829 -9864 -26811 -9819
rect -27270 -9891 -26811 -9864
rect -27378 -9954 -27360 -9891
rect -26829 -9918 -26811 -9891
rect -26667 -9918 -26649 -9819
rect -26370 -9828 -26352 -9792
rect -26361 -9855 -26352 -9828
rect -26370 -9864 -26352 -9855
rect -26370 -9909 -26352 -9891
rect -26829 -9954 -26811 -9945
rect -26667 -9954 -26649 -9945
rect -28170 -9990 -28152 -9981
rect -28044 -10107 -28026 -9981
rect -29016 -10134 -28026 -10107
rect -30285 -10170 -30123 -10152
rect -30069 -10170 -29871 -10152
rect -29808 -10170 -29763 -10152
rect -30330 -10296 -29961 -10278
rect -29781 -10368 -29763 -10170
rect -29520 -10350 -28188 -10332
rect -30177 -10548 -29736 -10530
rect -30177 -10638 -30159 -10548
rect -30330 -10656 -30123 -10638
rect -30069 -10656 -30060 -10638
rect -30042 -10656 -29871 -10638
rect -29808 -10656 -29781 -10638
rect -30879 -11187 -30366 -11169
rect -30330 -11295 -30312 -10656
rect -30042 -10809 -30024 -10656
rect -29754 -10809 -29736 -10548
rect -29475 -10692 -29457 -10674
rect -29475 -10782 -29457 -10746
rect -27900 -10773 -27882 -9981
rect -30285 -10827 -30123 -10809
rect -30069 -10827 -30024 -10809
rect -29907 -10827 -29871 -10809
rect -29808 -10827 -29736 -10809
rect -29691 -10809 -29511 -10782
rect -29466 -10809 -29457 -10782
rect -29385 -10800 -27882 -10773
rect -29475 -10818 -29457 -10809
rect -30285 -11169 -30267 -10827
rect -29475 -10863 -29457 -10845
rect -29997 -11007 -29961 -10980
rect -30186 -11025 -30123 -11007
rect -30069 -11025 -29871 -11007
rect -29808 -11025 -29763 -11007
rect -29997 -11169 -29961 -11124
rect -30240 -11187 -30123 -11169
rect -30069 -11187 -29871 -11169
rect -29808 -11187 -29790 -11169
rect -30330 -11313 -29961 -11295
rect -29781 -11403 -29763 -11025
rect -31077 -11421 -29763 -11403
rect -33840 -11538 -33822 -11511
rect -33678 -11538 -33660 -11511
rect -33840 -11646 -33822 -11583
rect -34011 -11664 -33822 -11646
rect -35379 -12078 -35361 -12069
rect -35379 -12123 -35361 -12105
rect -35676 -12132 -35658 -12123
rect -35838 -12168 -35820 -12159
rect -35676 -12168 -35658 -12159
rect -36171 -12231 -36153 -12195
rect -36423 -12258 -36153 -12231
rect -36423 -13095 -36405 -12258
rect -36171 -12267 -36153 -12258
rect -36171 -12312 -36153 -12294
rect -35379 -12393 -35361 -12276
rect -35838 -12429 -35820 -12402
rect -35676 -12429 -35658 -12402
rect -36162 -12465 -36144 -12447
rect -34011 -12420 -33993 -11664
rect -33840 -11682 -33822 -11664
rect -33678 -11682 -33660 -11583
rect -33381 -11592 -33363 -11556
rect -33372 -11619 -33363 -11592
rect -33291 -11610 -31257 -11583
rect -33381 -11628 -33363 -11619
rect -33381 -11673 -33363 -11655
rect -33840 -11718 -33822 -11709
rect -33678 -11763 -33660 -11709
rect -33165 -11718 -29349 -11682
rect -30177 -11844 -29736 -11826
rect -30177 -11934 -30159 -11844
rect -30330 -11952 -30123 -11934
rect -30069 -11952 -30060 -11934
rect -30042 -11952 -29871 -11934
rect -29808 -11952 -29781 -11934
rect -33381 -12366 -33363 -12249
rect -33840 -12402 -33822 -12375
rect -33678 -12402 -33660 -12375
rect -34137 -12438 -33993 -12420
rect -35838 -12519 -35820 -12474
rect -36162 -12555 -36144 -12519
rect -36369 -12582 -36144 -12555
rect -35838 -12573 -35820 -12537
rect -35676 -12546 -35658 -12474
rect -35379 -12483 -35361 -12447
rect -34137 -12474 -34119 -12438
rect -35370 -12510 -35361 -12483
rect -35289 -12501 -34119 -12474
rect -33840 -12510 -33822 -12447
rect -35379 -12519 -35361 -12510
rect -35703 -12564 -35658 -12546
rect -34011 -12528 -33822 -12510
rect -35379 -12564 -35361 -12546
rect -35703 -12573 -35685 -12564
rect -35676 -12573 -35658 -12564
rect -36369 -12699 -36351 -12582
rect -36162 -12591 -36144 -12582
rect -35838 -12609 -35820 -12600
rect -36162 -12636 -36144 -12618
rect -35703 -12699 -35685 -12600
rect -35676 -12609 -35658 -12600
rect -36369 -12717 -35685 -12699
rect -35982 -12924 -35964 -12717
rect -35379 -12807 -35361 -12690
rect -35838 -12843 -35820 -12816
rect -35676 -12843 -35658 -12816
rect -35838 -12924 -35820 -12888
rect -35982 -12942 -35820 -12924
rect -35838 -12987 -35820 -12942
rect -35676 -12960 -35658 -12888
rect -35379 -12897 -35361 -12861
rect -34011 -12888 -33993 -12528
rect -33840 -12546 -33822 -12528
rect -33678 -12546 -33660 -12447
rect -33381 -12456 -33363 -12420
rect -33372 -12483 -33363 -12456
rect -33381 -12492 -33363 -12483
rect -33381 -12537 -33363 -12519
rect -33840 -12582 -33822 -12573
rect -33678 -12618 -33660 -12573
rect -33318 -12582 -30411 -12555
rect -30330 -12591 -30312 -11952
rect -30042 -12105 -30024 -11952
rect -29754 -12105 -29736 -11844
rect -29475 -11988 -29457 -11970
rect -29475 -12078 -29457 -12042
rect -27774 -12069 -27756 -9981
rect -27639 -9990 -27621 -9981
rect -27378 -9990 -27360 -9981
rect -30285 -12123 -30123 -12105
rect -30069 -12123 -30024 -12105
rect -29907 -12123 -29871 -12105
rect -29808 -12123 -29736 -12105
rect -29691 -12105 -29511 -12078
rect -29466 -12105 -29457 -12078
rect -29385 -12096 -27756 -12069
rect -29475 -12114 -29457 -12105
rect -30285 -12465 -30267 -12123
rect -29475 -12159 -29457 -12141
rect -29997 -12303 -29961 -12276
rect -30141 -12321 -30123 -12303
rect -30069 -12321 -29871 -12303
rect -29808 -12321 -29763 -12303
rect -29997 -12465 -29961 -12420
rect -30285 -12483 -30123 -12465
rect -30069 -12483 -29871 -12465
rect -29808 -12483 -29763 -12465
rect -30330 -12609 -29961 -12591
rect -29781 -12681 -29763 -12483
rect -31356 -12699 -29763 -12681
rect -33381 -12861 -33363 -12744
rect -35370 -12924 -35361 -12897
rect -35289 -12915 -33993 -12888
rect -33840 -12897 -33822 -12870
rect -33678 -12897 -33660 -12870
rect -35379 -12933 -35361 -12924
rect -35721 -12978 -35658 -12960
rect -35379 -12978 -35361 -12960
rect -35721 -12987 -35703 -12978
rect -35676 -12987 -35658 -12978
rect -34011 -13005 -33993 -12915
rect -33840 -13005 -33822 -12942
rect -35838 -13023 -35820 -13014
rect -35721 -13095 -35703 -13014
rect -35676 -13023 -35658 -13014
rect -34011 -13023 -33822 -13005
rect -36423 -13113 -35703 -13095
rect -34011 -13428 -33993 -13023
rect -33840 -13041 -33822 -13023
rect -33678 -13041 -33660 -12942
rect -33381 -12951 -33363 -12915
rect -33372 -12978 -33363 -12951
rect -33381 -12987 -33363 -12978
rect -33381 -13032 -33363 -13014
rect -33840 -13077 -33822 -13068
rect -33678 -13113 -33660 -13068
rect -33381 -13275 -33363 -13158
rect -33840 -13311 -33822 -13284
rect -33678 -13311 -33660 -13284
rect -33840 -13428 -33822 -13356
rect -34011 -13446 -33822 -13428
rect -34011 -13950 -33993 -13446
rect -33840 -13455 -33822 -13446
rect -33678 -13455 -33660 -13356
rect -33381 -13365 -33363 -13329
rect -33372 -13392 -33363 -13365
rect -33381 -13401 -33363 -13392
rect -33381 -13446 -33363 -13428
rect -33840 -13491 -33822 -13482
rect -33678 -13554 -33660 -13482
rect -33381 -13806 -33363 -13689
rect -33840 -13842 -33822 -13815
rect -33678 -13842 -33660 -13815
rect -31410 -13815 -31392 -13698
rect -31869 -13851 -31851 -13824
rect -31707 -13851 -31689 -13824
rect -33840 -13950 -33822 -13887
rect -34011 -13968 -33822 -13950
rect -34011 -14445 -33993 -13968
rect -33840 -13986 -33822 -13968
rect -33678 -13986 -33660 -13887
rect -33381 -13896 -33363 -13860
rect -33372 -13923 -33363 -13896
rect -33381 -13932 -33363 -13923
rect -33381 -13977 -33363 -13959
rect -31869 -13995 -31851 -13896
rect -31707 -13995 -31689 -13896
rect -31410 -13905 -31392 -13869
rect -31401 -13932 -31392 -13905
rect -31410 -13941 -31392 -13932
rect -31410 -13986 -31392 -13968
rect -33840 -14022 -33822 -14013
rect -33678 -14067 -33660 -14013
rect -31869 -14076 -31851 -14022
rect -31707 -14076 -31689 -14022
rect -33381 -14301 -33363 -14184
rect -31410 -14292 -31392 -14175
rect -33840 -14337 -33822 -14310
rect -33678 -14337 -33660 -14310
rect -31869 -14328 -31851 -14301
rect -31707 -14328 -31689 -14301
rect -33840 -14445 -33822 -14382
rect -34011 -14463 -33822 -14445
rect -34011 -14940 -33993 -14463
rect -33840 -14481 -33822 -14463
rect -33678 -14481 -33660 -14382
rect -33381 -14391 -33363 -14355
rect -33372 -14418 -33363 -14391
rect -33381 -14427 -33363 -14418
rect -33381 -14472 -33363 -14454
rect -31869 -14472 -31851 -14373
rect -31707 -14472 -31689 -14373
rect -31410 -14382 -31392 -14346
rect -31401 -14409 -31392 -14382
rect -31410 -14418 -31392 -14409
rect -31410 -14463 -31392 -14445
rect -33840 -14517 -33822 -14508
rect -33678 -14562 -33660 -14508
rect -31869 -14544 -31851 -14499
rect -31707 -14544 -31689 -14499
rect -33381 -14796 -33363 -14679
rect -31410 -14688 -31392 -14571
rect -31869 -14724 -31851 -14697
rect -31707 -14724 -31689 -14697
rect -33840 -14832 -33822 -14805
rect -33678 -14832 -33660 -14805
rect -33840 -14940 -33822 -14877
rect -34011 -14958 -33822 -14940
rect -34011 -15363 -33993 -14958
rect -33840 -14976 -33822 -14958
rect -33678 -14976 -33660 -14877
rect -33381 -14886 -33363 -14850
rect -31869 -14868 -31851 -14769
rect -31707 -14868 -31689 -14769
rect -31410 -14778 -31392 -14742
rect -31401 -14805 -31392 -14778
rect -31410 -14814 -31392 -14805
rect -31410 -14859 -31392 -14841
rect -33372 -14913 -33363 -14886
rect -33381 -14922 -33363 -14913
rect -31869 -14940 -31851 -14895
rect -33381 -14967 -33363 -14949
rect -31707 -14940 -31689 -14895
rect -33840 -15012 -33822 -15003
rect -33678 -15048 -33660 -15003
rect -33381 -15210 -33363 -15093
rect -31410 -15156 -31392 -15039
rect -31869 -15192 -31851 -15165
rect -31707 -15192 -31689 -15165
rect -33840 -15246 -33822 -15219
rect -33678 -15246 -33660 -15219
rect -33840 -15363 -33822 -15291
rect -34011 -15381 -33822 -15363
rect -34011 -15885 -33993 -15381
rect -33840 -15390 -33822 -15381
rect -33678 -15390 -33660 -15291
rect -33381 -15300 -33363 -15264
rect -33372 -15327 -33363 -15300
rect -33381 -15336 -33363 -15327
rect -31869 -15336 -31851 -15237
rect -31707 -15336 -31689 -15237
rect -31410 -15246 -31392 -15210
rect -31401 -15273 -31392 -15246
rect -31410 -15282 -31392 -15273
rect -31410 -15327 -31392 -15309
rect -33381 -15381 -33363 -15363
rect -31869 -15417 -31851 -15363
rect -33840 -15426 -33822 -15417
rect -33678 -15471 -33660 -15417
rect -31707 -15417 -31689 -15363
rect -33381 -15741 -33363 -15624
rect -33840 -15777 -33822 -15750
rect -33678 -15777 -33660 -15750
rect -33840 -15885 -33822 -15822
rect -34011 -15903 -33822 -15885
rect -33840 -15921 -33822 -15903
rect -33678 -15921 -33660 -15822
rect -33381 -15831 -33363 -15795
rect -33372 -15858 -33363 -15831
rect -33381 -15867 -33363 -15858
rect -33381 -15912 -33363 -15894
rect -33840 -15957 -33822 -15948
rect -33678 -16002 -33660 -15948
<< polycontact >>
rect -30852 9882 -30834 9900
rect -30087 10170 -30051 10188
rect -30357 9945 -30321 9981
rect -30537 9828 -30519 9855
rect -30348 9765 -30330 9801
rect -30357 9630 -30321 9666
rect -29970 9864 -29952 9882
rect -29277 10170 -29241 10188
rect -29547 9945 -29511 9981
rect -29718 9819 -29691 9846
rect -29538 9738 -29520 9765
rect -29547 9630 -29511 9666
rect -29088 9855 -29070 9882
rect -28395 10152 -28359 10197
rect -28665 9945 -28629 9981
rect -28836 9819 -28809 9846
rect -28656 9765 -28638 9792
rect -28665 9630 -28629 9666
rect -28521 9639 -28494 9657
rect -29538 9477 -29511 9495
rect -29610 9432 -29592 9450
rect -29889 9261 -29862 9288
rect -29808 9270 -29772 9297
rect -28989 9549 -28971 9567
rect -28863 9324 -28836 9351
rect -28782 9333 -28746 9360
rect -28989 9198 -28971 9216
rect -29529 9171 -29511 9189
rect -29610 9009 -29592 9027
rect -29439 8874 -29430 8892
rect -30852 7785 -30834 7803
rect -30087 8073 -30051 8091
rect -30357 7848 -30321 7884
rect -30546 7731 -30528 7758
rect -30348 7677 -30330 7704
rect -30357 7533 -30321 7569
rect -29970 7767 -29952 7785
rect -29277 8073 -29241 8091
rect -29547 7848 -29511 7884
rect -29718 7722 -29691 7749
rect -29538 7641 -29520 7668
rect -29547 7533 -29511 7569
rect -29088 7758 -29070 7785
rect -28395 8055 -28359 8100
rect -28665 7848 -28629 7884
rect -28836 7722 -28809 7749
rect -28656 7677 -28638 7704
rect -28665 7533 -28629 7569
rect -28521 7551 -28485 7569
rect -29538 7380 -29511 7398
rect -29610 7335 -29592 7353
rect -29889 7164 -29862 7191
rect -29808 7173 -29772 7200
rect -28989 7452 -28971 7470
rect -28863 7227 -28836 7254
rect -28782 7236 -28746 7263
rect -28989 7101 -28971 7119
rect -29529 7074 -29511 7092
rect -29610 6912 -29592 6930
rect -29439 6777 -29430 6795
rect -30852 5670 -30834 5688
rect -30087 5958 -30051 5976
rect -30357 5733 -30321 5769
rect -30546 5616 -30528 5643
rect -30348 5553 -30330 5589
rect -30357 5418 -30321 5454
rect -29970 5652 -29952 5670
rect -29277 5958 -29241 5976
rect -29547 5733 -29511 5769
rect -29718 5607 -29691 5634
rect -29538 5526 -29511 5553
rect -29547 5418 -29511 5454
rect -29088 5643 -29070 5670
rect -28395 5940 -28359 5985
rect -28665 5733 -28629 5769
rect -28836 5607 -28809 5634
rect -28656 5562 -28638 5580
rect -28665 5418 -28629 5454
rect -29538 5265 -29511 5283
rect -29610 5220 -29592 5238
rect -29889 5049 -29862 5076
rect -29808 5058 -29772 5085
rect -28989 5337 -28971 5355
rect -28863 5112 -28836 5139
rect -28782 5121 -28746 5148
rect -28989 4986 -28971 5004
rect -29529 4959 -29511 4977
rect -29610 4797 -29592 4815
rect -27792 6777 -27765 6795
rect -29439 4662 -29430 4680
rect -29403 4662 -29367 4680
rect -30726 3807 -30708 3825
rect -30726 3762 -30708 3789
rect -30087 4023 -30051 4041
rect -30357 3798 -30321 3834
rect -30528 3726 -30510 3744
rect -30348 3627 -30330 3654
rect -30357 3483 -30321 3519
rect -29970 3717 -29952 3735
rect -29277 4023 -29241 4041
rect -29547 3798 -29511 3834
rect -29718 3672 -29691 3699
rect -29538 3591 -29511 3618
rect -29547 3483 -29511 3519
rect -29088 3708 -29070 3735
rect -28395 4005 -28359 4050
rect -28665 3798 -28629 3834
rect -28836 3672 -28809 3699
rect -28656 3627 -28638 3645
rect -28665 3483 -28629 3519
rect -29538 3330 -29511 3348
rect -29610 3285 -29592 3303
rect -29889 3114 -29862 3141
rect -29808 3123 -29772 3150
rect -28989 3402 -28971 3420
rect -28350 3348 -28332 3411
rect -28863 3177 -28836 3204
rect -28782 3186 -28746 3213
rect -28989 3051 -28971 3069
rect -29529 3024 -29511 3042
rect -29610 2862 -29592 2880
rect -29439 2727 -29430 2745
rect -36801 1035 -36783 1152
rect -30744 -99 -30699 -81
rect -30366 -99 -30339 -81
rect -29718 270 -29691 306
rect -29511 279 -29466 306
rect -29448 189 -29421 207
rect -29997 108 -29961 144
rect -30168 63 -30141 81
rect -29988 -27 -29970 -9
rect -30285 -99 -30249 -81
rect -29997 -207 -29961 -171
rect -28431 135 -28404 153
rect -29124 -27 -29097 0
rect -29043 -18 -29016 9
rect -28287 9 -28260 36
rect -27045 18 -27018 45
rect -29151 -117 -29124 -99
rect -33417 -405 -33390 -378
rect -33696 -585 -33678 -549
rect -33696 -747 -33678 -702
rect -33417 -900 -33390 -873
rect -30969 -1053 -30942 -1017
rect -30915 -1044 -30879 -1026
rect -30366 -1044 -30339 -1026
rect -34209 -1179 -34200 -1161
rect -34164 -1179 -34119 -1161
rect -36801 -1413 -36783 -1341
rect -33417 -1314 -33390 -1287
rect -33696 -1494 -33678 -1458
rect -33417 -1845 -33390 -1818
rect -33696 -2052 -33678 -1989
rect -33417 -2412 -33390 -2385
rect -33696 -2601 -33678 -2547
rect -33417 -2907 -33390 -2880
rect -33696 -3078 -33678 -3051
rect -33417 -3321 -33390 -3294
rect -33696 -3519 -33678 -3474
rect -31023 -3744 -30987 -3726
rect -33417 -3852 -33390 -3825
rect -33696 -4041 -33678 -3987
rect -31284 -6723 -31266 -6687
rect -29718 -675 -29691 -639
rect -29511 -666 -29466 -639
rect -27882 -576 -27864 -522
rect -29475 -756 -29457 -738
rect -29997 -837 -29961 -801
rect -30168 -882 -30132 -864
rect -29142 -837 -29115 -810
rect -29061 -828 -29016 -801
rect -28359 -801 -28332 -774
rect -28278 -792 -28242 -765
rect -27531 -801 -27504 -774
rect -27090 -819 -27072 -801
rect -26919 -810 -26892 -792
rect -26820 -810 -26802 -792
rect -26694 -837 -26685 -819
rect -29169 -927 -29124 -909
rect -29988 -972 -29970 -954
rect -30285 -1044 -30249 -1026
rect -29997 -1152 -29961 -1116
rect -30924 -2061 -30888 -2043
rect -30366 -2061 -30339 -2043
rect -28656 -1629 -28629 -1602
rect -27855 -1611 -27828 -1584
rect -29718 -1692 -29691 -1656
rect -29511 -1683 -29466 -1656
rect -29160 -1683 -29133 -1656
rect -28521 -1647 -28494 -1620
rect -28377 -1647 -28350 -1620
rect -28251 -1647 -28224 -1620
rect -28116 -1647 -28089 -1620
rect -29457 -1773 -29421 -1755
rect -29178 -1773 -29142 -1755
rect -29997 -1854 -29961 -1818
rect -29943 -1980 -29925 -1962
rect -29988 -2034 -29970 -2007
rect -30285 -2061 -30249 -2043
rect -29997 -2169 -29961 -2133
rect -29916 -2196 -29898 -2169
rect -30771 -2340 -30735 -2322
rect -28809 -2925 -28782 -2898
rect -28008 -2907 -27981 -2880
rect -29718 -2988 -29691 -2952
rect -29511 -2979 -29466 -2952
rect -29214 -2979 -29187 -2952
rect -28674 -2943 -28647 -2916
rect -28530 -2943 -28503 -2916
rect -28404 -2943 -28377 -2916
rect -28269 -2943 -28242 -2916
rect -29997 -3150 -29961 -3114
rect -29610 -3240 -29583 -3195
rect -29943 -3276 -29925 -3249
rect -29988 -3321 -29970 -3303
rect -29997 -3465 -29961 -3429
rect -29610 -3915 -29583 -3861
rect -29718 -4059 -29691 -4023
rect -29511 -4050 -29466 -4023
rect -29448 -4140 -29421 -4122
rect -29997 -4221 -29961 -4185
rect -29988 -4356 -29970 -4338
rect -29997 -4536 -29961 -4500
rect -29124 -4356 -29097 -4329
rect -29043 -4347 -29016 -4320
rect -28287 -4320 -28260 -4293
rect -27045 -4311 -27018 -4284
rect -29151 -4446 -29124 -4428
rect -30852 -4680 -30780 -4662
rect -30960 -5409 -30942 -5373
rect -29718 -5004 -29691 -4968
rect -29511 -4995 -29466 -4968
rect -27882 -4905 -27864 -4851
rect -29475 -5085 -29457 -5067
rect -29997 -5166 -29961 -5130
rect -29142 -5166 -29115 -5139
rect -29061 -5157 -29016 -5130
rect -28359 -5130 -28332 -5103
rect -28278 -5121 -28242 -5094
rect -27531 -5130 -27504 -5103
rect -27090 -5148 -27072 -5130
rect -26919 -5139 -26892 -5121
rect -26820 -5139 -26802 -5121
rect -26694 -5166 -26685 -5148
rect -29169 -5256 -29124 -5238
rect -29988 -5301 -29970 -5283
rect -30240 -5373 -30213 -5355
rect -29997 -5481 -29961 -5445
rect -30240 -5526 -30213 -5508
rect -31131 -5688 -31086 -5670
rect -28656 -5958 -28629 -5931
rect -27855 -5940 -27828 -5913
rect -29718 -6021 -29691 -5985
rect -29511 -6012 -29466 -5985
rect -29160 -6012 -29133 -5985
rect -28521 -5976 -28494 -5949
rect -28377 -5976 -28350 -5949
rect -28251 -5976 -28224 -5949
rect -28116 -5976 -28089 -5949
rect -29457 -6102 -29421 -6084
rect -29178 -6102 -29142 -6084
rect -29997 -6183 -29961 -6147
rect -29943 -6309 -29925 -6291
rect -29988 -6363 -29970 -6336
rect -30240 -6390 -30222 -6372
rect -29997 -6498 -29961 -6462
rect -29943 -6534 -29925 -6498
rect -31167 -7947 -31149 -7902
rect -31077 -6642 -31050 -6606
rect -33399 -8262 -33372 -8235
rect -33336 -8253 -33291 -8226
rect -33687 -8433 -33651 -8406
rect -33399 -8757 -33372 -8730
rect -33327 -8748 -33291 -8721
rect -31545 -8748 -31500 -8721
rect -33678 -8928 -33660 -8901
rect -33399 -9171 -33372 -9144
rect -33318 -9162 -33291 -9135
rect -31437 -9153 -31419 -9126
rect -33678 -9351 -33660 -9315
rect -31284 -9414 -31266 -9387
rect -33399 -9702 -33372 -9675
rect -33327 -9693 -33291 -9666
rect -31437 -9693 -31392 -9666
rect -33678 -9891 -33651 -9855
rect -33399 -10179 -33372 -10152
rect -33327 -10170 -33291 -10143
rect -33687 -10359 -33651 -10332
rect -31455 -10467 -31383 -10449
rect -35847 -11637 -35820 -11619
rect -35397 -11601 -35370 -11574
rect -35325 -11592 -35289 -11565
rect -35694 -11655 -35658 -11637
rect -35397 -12069 -35370 -12042
rect -35334 -12060 -35289 -12033
rect -33399 -10674 -33372 -10647
rect -33327 -10665 -33291 -10638
rect -31518 -10665 -31473 -10638
rect -33678 -10854 -33660 -10818
rect -30879 -7065 -30861 -7020
rect -30960 -10368 -30942 -10341
rect -30960 -10665 -30942 -10602
rect -33399 -11088 -33372 -11061
rect -33327 -11079 -33291 -11052
rect -33678 -11259 -33660 -11232
rect -29340 -7137 -29322 -7065
rect -29718 -7317 -29691 -7281
rect -29511 -7308 -29466 -7281
rect -29997 -7479 -29961 -7443
rect -29943 -7605 -29925 -7578
rect -29988 -7650 -29970 -7632
rect -29997 -7794 -29961 -7758
rect -28809 -7254 -28782 -7227
rect -28008 -7236 -27981 -7209
rect -29214 -7308 -29187 -7281
rect -28674 -7272 -28647 -7245
rect -28530 -7272 -28503 -7245
rect -28404 -7272 -28377 -7245
rect -28269 -7272 -28242 -7245
rect -29340 -8721 -29322 -8631
rect -29718 -8856 -29691 -8820
rect -29511 -8847 -29466 -8820
rect -29412 -8838 -29385 -8811
rect -29997 -9018 -29961 -8982
rect -30186 -9063 -30168 -9045
rect -29997 -9333 -29961 -9297
rect -29781 -9450 -29763 -9432
rect -29718 -9801 -29691 -9765
rect -29511 -9792 -29466 -9765
rect -29412 -9783 -29385 -9756
rect -29997 -9963 -29961 -9927
rect -30186 -10008 -30168 -9990
rect -27387 -9891 -27360 -9864
rect -27324 -9891 -27270 -9864
rect -26388 -9855 -26361 -9828
rect -29997 -10278 -29961 -10242
rect -29556 -10350 -29520 -10332
rect -28188 -10350 -28170 -10314
rect -29781 -10404 -29763 -10368
rect -30366 -11187 -30339 -11169
rect -29718 -10818 -29691 -10782
rect -29511 -10809 -29466 -10782
rect -29412 -10800 -29385 -10773
rect -29997 -10980 -29961 -10944
rect -30285 -11187 -30240 -11169
rect -29997 -11295 -29961 -11259
rect -35676 -12123 -35658 -12105
rect -33399 -11619 -33372 -11592
rect -33336 -11610 -33291 -11583
rect -31257 -11610 -31203 -11583
rect -33210 -11718 -33165 -11682
rect -29349 -11718 -29313 -11673
rect -33678 -11826 -33660 -11763
rect -35838 -12537 -35820 -12519
rect -35397 -12510 -35370 -12483
rect -35334 -12501 -35289 -12474
rect -33399 -12483 -33372 -12456
rect -33381 -12582 -33318 -12555
rect -30411 -12600 -30375 -12546
rect -29718 -12114 -29691 -12078
rect -29511 -12105 -29466 -12078
rect -29412 -12096 -29385 -12069
rect -29997 -12276 -29961 -12240
rect -30168 -12321 -30141 -12303
rect -29997 -12591 -29961 -12555
rect -33678 -12645 -33660 -12618
rect -31374 -12699 -31356 -12681
rect -35397 -12924 -35370 -12897
rect -35334 -12915 -35289 -12888
rect -33399 -12978 -33372 -12951
rect -33678 -13131 -33660 -13113
rect -33399 -13392 -33372 -13365
rect -33678 -13590 -33660 -13554
rect -33399 -13923 -33372 -13896
rect -31428 -13932 -31401 -13905
rect -33687 -14094 -33651 -14067
rect -31869 -14112 -31851 -14076
rect -31707 -14103 -31689 -14076
rect -33399 -14418 -33372 -14391
rect -31428 -14409 -31401 -14382
rect -33678 -14598 -33660 -14562
rect -31869 -14571 -31851 -14544
rect -31707 -14580 -31689 -14544
rect -31428 -14805 -31401 -14778
rect -33399 -14913 -33372 -14886
rect -31869 -14967 -31851 -14940
rect -31707 -15003 -31689 -14940
rect -33678 -15075 -33660 -15048
rect -33399 -15327 -33372 -15300
rect -31428 -15273 -31401 -15246
rect -31869 -15471 -31851 -15417
rect -33678 -15516 -33660 -15471
rect -31707 -15480 -31689 -15417
rect -33399 -15858 -33372 -15831
rect -33678 -16047 -33660 -16002
<< metal1 >>
rect -29574 10467 -29538 10485
rect -30438 10296 -30222 10332
rect -30186 10296 -30006 10332
rect -29628 10296 -29412 10332
rect -29376 10296 -29196 10332
rect -28746 10296 -28530 10332
rect -28494 10296 -28314 10332
rect -30438 10224 -30222 10260
rect -30186 10224 -30051 10260
rect -30087 10188 -30051 10224
rect -30600 10125 -30474 10161
rect -30438 10125 -30222 10161
rect -30600 10026 -30564 10125
rect -30087 10089 -30051 10170
rect -30438 10053 -30222 10089
rect -30186 10053 -30051 10089
rect -30042 10026 -30006 10296
rect -29628 10224 -29412 10260
rect -29376 10224 -29241 10260
rect -29277 10188 -29241 10224
rect -30600 9990 -30375 10026
rect -30600 9936 -30474 9972
rect -30834 9882 -30798 9900
rect -30600 9873 -30564 9900
rect -30753 9855 -30564 9873
rect -30753 9153 -30735 9855
rect -30600 9846 -30564 9855
rect -30411 9891 -30375 9990
rect -30357 9990 -30006 10026
rect -29790 10125 -29664 10161
rect -29628 10125 -29412 10161
rect -29790 10026 -29754 10125
rect -29277 10089 -29241 10170
rect -29628 10053 -29412 10089
rect -29376 10053 -29241 10089
rect -29232 10026 -29196 10296
rect -28746 10224 -28530 10260
rect -28494 10224 -28359 10260
rect -28395 10197 -28359 10224
rect -29790 9990 -29565 10026
rect -30357 9981 -30321 9990
rect -30186 9936 -30069 9972
rect -30537 9855 -30519 9873
rect -30438 9855 -30222 9891
rect -30105 9873 -30069 9900
rect -29790 9936 -29664 9972
rect -30105 9855 -29979 9873
rect -29952 9864 -29898 9882
rect -30105 9846 -30069 9855
rect -30600 9774 -30474 9810
rect -30186 9774 -30069 9810
rect -30438 9693 -30222 9729
rect -30357 9666 -30321 9693
rect -29997 9405 -29979 9855
rect -29790 9846 -29754 9900
rect -29601 9891 -29565 9990
rect -29547 9990 -29196 10026
rect -28908 10125 -28782 10161
rect -28746 10125 -28530 10161
rect -28908 10026 -28872 10125
rect -28395 10089 -28359 10152
rect -28746 10053 -28530 10089
rect -28494 10053 -28359 10089
rect -28350 10026 -28314 10296
rect -28908 9990 -28683 10026
rect -29547 9981 -29511 9990
rect -29376 9936 -29259 9972
rect -29628 9855 -29412 9891
rect -29295 9882 -29259 9900
rect -28908 9936 -28782 9972
rect -28908 9882 -28872 9900
rect -28719 9891 -28683 9990
rect -28665 9990 -28314 10026
rect -28665 9981 -28629 9990
rect -28494 9936 -28377 9972
rect -29295 9864 -29178 9882
rect -29718 9846 -29700 9855
rect -29295 9846 -29259 9864
rect -29790 9774 -29664 9810
rect -29718 9495 -29700 9774
rect -29376 9774 -29259 9810
rect -29628 9693 -29412 9729
rect -29547 9666 -29511 9693
rect -29718 9477 -29538 9495
rect -29196 9468 -29178 9864
rect -29070 9855 -29043 9882
rect -28917 9864 -28872 9882
rect -28908 9846 -28872 9864
rect -28746 9855 -28530 9891
rect -28413 9882 -28377 9900
rect -28413 9864 -28386 9882
rect -28836 9846 -28809 9855
rect -28413 9846 -28377 9864
rect -28908 9774 -28782 9810
rect -28881 9567 -28863 9774
rect -28494 9774 -28377 9810
rect -28746 9693 -28530 9729
rect -28665 9666 -28629 9693
rect -28530 9639 -28521 9657
rect -28971 9549 -28863 9567
rect -28350 9513 -28332 9864
rect -28881 9495 -28332 9513
rect -28881 9468 -28854 9495
rect -29331 9450 -28854 9468
rect -29907 9432 -29610 9450
rect -29592 9432 -29313 9450
rect -29907 9405 -29880 9432
rect -30357 9387 -29880 9405
rect -30357 9333 -30339 9387
rect -30204 9333 -30186 9387
rect -29907 9378 -29880 9387
rect -29331 9396 -29313 9432
rect -29178 9396 -29160 9450
rect -28881 9441 -28854 9450
rect -30303 9252 -30285 9306
rect -30141 9252 -30123 9315
rect -29979 9261 -29889 9288
rect -29979 9252 -29961 9261
rect -30303 9234 -29961 9252
rect -29835 9252 -29808 9342
rect -29277 9315 -29259 9369
rect -29115 9315 -29097 9378
rect -28953 9324 -28863 9351
rect -28953 9315 -28935 9324
rect -29277 9297 -28935 9315
rect -28809 9315 -28782 9405
rect -29115 9261 -29097 9297
rect -30141 9198 -30123 9234
rect -28881 9252 -28854 9279
rect -29907 9189 -29880 9216
rect -29331 9216 -29313 9234
rect -28881 9234 -28782 9252
rect -28881 9216 -28845 9234
rect -29331 9198 -28989 9216
rect -28971 9198 -28845 9216
rect -29331 9189 -29313 9198
rect -30357 9153 -30339 9171
rect -29907 9171 -29529 9189
rect -29511 9171 -29313 9189
rect -29907 9153 -29871 9171
rect -31104 9135 -29871 9153
rect -31104 7056 -31086 9135
rect -29889 8802 -29871 9135
rect -29691 9009 -29610 9027
rect -29592 9009 -29421 9027
rect -29691 8973 -29673 9009
rect -29466 8973 -29448 9009
rect -29538 8892 -29520 8946
rect -29412 8892 -29394 8946
rect -29628 8874 -29439 8892
rect -29412 8874 -29367 8892
rect -29628 8847 -29610 8874
rect -29538 8847 -29520 8874
rect -29412 8847 -29394 8874
rect -29682 8802 -29664 8829
rect -29592 8802 -29574 8829
rect -29466 8802 -29448 8829
rect -29889 8784 -29448 8802
rect -29547 8370 -29538 8388
rect -30438 8199 -30222 8235
rect -30186 8199 -30006 8235
rect -29628 8199 -29412 8235
rect -29376 8199 -29196 8235
rect -28746 8199 -28530 8235
rect -28494 8199 -28314 8235
rect -30438 8127 -30222 8163
rect -30186 8127 -30051 8163
rect -30087 8091 -30051 8127
rect -30600 8028 -30474 8064
rect -30438 8028 -30222 8064
rect -30600 7929 -30564 8028
rect -30087 7992 -30051 8073
rect -30438 7956 -30222 7992
rect -30186 7956 -30051 7992
rect -30042 7929 -30006 8199
rect -29628 8127 -29412 8163
rect -29376 8127 -29241 8163
rect -29277 8091 -29241 8127
rect -30600 7893 -30375 7929
rect -30600 7839 -30474 7875
rect -30834 7785 -30816 7803
rect -30600 7776 -30564 7803
rect -30411 7794 -30375 7893
rect -30357 7893 -30006 7929
rect -29790 8028 -29664 8064
rect -29628 8028 -29412 8064
rect -29790 7929 -29754 8028
rect -29277 7992 -29241 8073
rect -29628 7956 -29412 7992
rect -29376 7956 -29241 7992
rect -29232 7929 -29196 8199
rect -28746 8127 -28530 8163
rect -28494 8127 -28359 8163
rect -28395 8100 -28359 8127
rect -29790 7893 -29565 7929
rect -30357 7884 -30321 7893
rect -30186 7839 -30069 7875
rect -30753 7758 -30564 7776
rect -30753 7056 -30735 7758
rect -30600 7749 -30564 7758
rect -30546 7758 -30528 7785
rect -30438 7758 -30222 7794
rect -30105 7776 -30069 7803
rect -29790 7839 -29664 7875
rect -30105 7758 -29979 7776
rect -29952 7767 -29898 7785
rect -30105 7749 -30069 7758
rect -30600 7677 -30474 7713
rect -30186 7677 -30069 7713
rect -30438 7596 -30222 7632
rect -30357 7569 -30321 7596
rect -29997 7308 -29979 7758
rect -29790 7749 -29754 7803
rect -29601 7794 -29565 7893
rect -29547 7893 -29196 7929
rect -28908 8028 -28782 8064
rect -28746 8028 -28530 8064
rect -28908 7929 -28872 8028
rect -28395 7992 -28359 8055
rect -28746 7956 -28530 7992
rect -28494 7956 -28359 7992
rect -28350 7929 -28314 8199
rect -28908 7893 -28683 7929
rect -29547 7884 -29511 7893
rect -29376 7839 -29259 7875
rect -29628 7758 -29412 7794
rect -29295 7785 -29259 7803
rect -28908 7839 -28782 7875
rect -28908 7785 -28872 7803
rect -28719 7794 -28683 7893
rect -28665 7893 -28314 7929
rect -28665 7884 -28629 7893
rect -28494 7839 -28377 7875
rect -29295 7767 -29178 7785
rect -29718 7749 -29700 7758
rect -29295 7749 -29259 7767
rect -29790 7677 -29664 7713
rect -29718 7398 -29700 7677
rect -29376 7677 -29259 7713
rect -29628 7596 -29412 7632
rect -29547 7569 -29511 7596
rect -29718 7380 -29538 7398
rect -29196 7371 -29178 7767
rect -29070 7758 -29043 7785
rect -28917 7767 -28872 7785
rect -28908 7749 -28872 7767
rect -28746 7758 -28530 7794
rect -28413 7785 -28377 7803
rect -28413 7767 -28386 7785
rect -28341 7767 -28332 7785
rect -28836 7749 -28809 7758
rect -28413 7749 -28377 7767
rect -28908 7677 -28782 7713
rect -28494 7677 -28377 7713
rect -28881 7470 -28863 7677
rect -28656 7668 -28638 7677
rect -28746 7596 -28530 7632
rect -28665 7569 -28629 7596
rect -28539 7551 -28521 7569
rect -28971 7452 -28863 7470
rect -28350 7416 -28332 7767
rect -28881 7398 -28332 7416
rect -28881 7371 -28854 7398
rect -29331 7353 -28854 7371
rect -29907 7335 -29610 7353
rect -29592 7335 -29313 7353
rect -29907 7308 -29880 7335
rect -30357 7290 -29880 7308
rect -30357 7236 -30339 7290
rect -30204 7236 -30186 7290
rect -29907 7281 -29880 7290
rect -29331 7299 -29313 7335
rect -29178 7299 -29160 7353
rect -28881 7344 -28854 7353
rect -30303 7155 -30285 7209
rect -30141 7155 -30123 7218
rect -29979 7164 -29889 7191
rect -29979 7155 -29961 7164
rect -30303 7137 -29961 7155
rect -29835 7155 -29808 7245
rect -29277 7218 -29259 7272
rect -29115 7218 -29097 7281
rect -28953 7227 -28863 7254
rect -28953 7218 -28935 7227
rect -29277 7200 -28935 7218
rect -28809 7218 -28782 7308
rect -29115 7164 -29097 7200
rect -30141 7101 -30123 7137
rect -28881 7155 -28854 7182
rect -29907 7092 -29880 7119
rect -29331 7119 -29313 7137
rect -28881 7137 -28782 7155
rect -28881 7119 -28845 7137
rect -29331 7101 -28989 7119
rect -28971 7101 -28845 7119
rect -29331 7092 -29313 7101
rect -30357 7056 -30339 7074
rect -29907 7074 -29529 7092
rect -29511 7074 -29313 7092
rect -29907 7056 -29871 7074
rect -31104 7038 -29871 7056
rect -31104 4941 -31086 7038
rect -29889 6705 -29871 7038
rect -29691 6912 -29610 6930
rect -29592 6912 -29421 6930
rect -29691 6876 -29673 6912
rect -29466 6876 -29448 6912
rect -29538 6795 -29520 6849
rect -29412 6795 -29394 6849
rect -29628 6777 -29439 6795
rect -29412 6777 -27792 6795
rect -29628 6750 -29610 6777
rect -29538 6750 -29520 6777
rect -29412 6750 -29394 6777
rect -29682 6705 -29664 6732
rect -29592 6705 -29574 6732
rect -29466 6705 -29448 6732
rect -29889 6687 -29448 6705
rect -29565 6228 -29538 6264
rect -30438 6084 -30222 6120
rect -30186 6084 -30006 6120
rect -29628 6084 -29412 6120
rect -29376 6084 -29196 6120
rect -28746 6084 -28530 6120
rect -28494 6084 -28314 6120
rect -30438 6012 -30222 6048
rect -30186 6012 -30051 6048
rect -30087 5976 -30051 6012
rect -30600 5913 -30474 5949
rect -30438 5913 -30222 5949
rect -30600 5814 -30564 5913
rect -30087 5877 -30051 5958
rect -30438 5841 -30222 5877
rect -30186 5841 -30051 5877
rect -30042 5814 -30006 6084
rect -29628 6012 -29412 6048
rect -29376 6012 -29241 6048
rect -29277 5976 -29241 6012
rect -30600 5778 -30375 5814
rect -30600 5724 -30474 5760
rect -30834 5670 -30816 5688
rect -30600 5661 -30564 5688
rect -30411 5679 -30375 5778
rect -30357 5778 -30006 5814
rect -29790 5913 -29664 5949
rect -29628 5913 -29412 5949
rect -29790 5814 -29754 5913
rect -29277 5877 -29241 5958
rect -29628 5841 -29412 5877
rect -29376 5841 -29241 5877
rect -29232 5814 -29196 6084
rect -28746 6012 -28530 6048
rect -28494 6012 -28359 6048
rect -28395 5985 -28359 6012
rect -29790 5778 -29565 5814
rect -30357 5769 -30321 5778
rect -30186 5724 -30069 5760
rect -30753 5643 -30564 5661
rect -30753 4941 -30735 5643
rect -30600 5634 -30564 5643
rect -30546 5643 -30528 5670
rect -30438 5643 -30222 5679
rect -30105 5661 -30069 5688
rect -29790 5724 -29664 5760
rect -30105 5643 -29979 5661
rect -29952 5652 -29898 5670
rect -30105 5634 -30069 5643
rect -30600 5562 -30474 5598
rect -30186 5562 -30069 5598
rect -30438 5481 -30222 5517
rect -30357 5454 -30321 5481
rect -29997 5193 -29979 5643
rect -29790 5634 -29754 5688
rect -29601 5679 -29565 5778
rect -29547 5778 -29196 5814
rect -28908 5913 -28782 5949
rect -28746 5913 -28530 5949
rect -28908 5814 -28872 5913
rect -28395 5877 -28359 5940
rect -28746 5841 -28530 5877
rect -28494 5841 -28359 5877
rect -28350 5814 -28314 6084
rect -28908 5778 -28683 5814
rect -29547 5769 -29511 5778
rect -29376 5724 -29259 5760
rect -29628 5643 -29412 5679
rect -29295 5670 -29259 5688
rect -28908 5724 -28782 5760
rect -28908 5670 -28872 5688
rect -28719 5679 -28683 5778
rect -28665 5778 -28314 5814
rect -28665 5769 -28629 5778
rect -28494 5724 -28377 5760
rect -29295 5652 -29178 5670
rect -29718 5634 -29700 5643
rect -29295 5634 -29259 5652
rect -29790 5562 -29664 5598
rect -29718 5283 -29700 5562
rect -29376 5562 -29259 5598
rect -29628 5481 -29412 5517
rect -29547 5454 -29511 5481
rect -29718 5265 -29538 5283
rect -29196 5256 -29178 5652
rect -29070 5643 -29043 5670
rect -28917 5652 -28872 5670
rect -28908 5634 -28872 5652
rect -28746 5643 -28530 5679
rect -28413 5670 -28377 5688
rect -28413 5652 -28368 5670
rect -28836 5634 -28809 5643
rect -28413 5634 -28377 5652
rect -28908 5562 -28782 5598
rect -28494 5562 -28377 5598
rect -28881 5355 -28863 5562
rect -28746 5481 -28530 5517
rect -28665 5454 -28629 5481
rect -28971 5337 -28863 5355
rect -28350 5301 -28332 5652
rect -28881 5283 -28332 5301
rect -28881 5256 -28854 5283
rect -29331 5238 -28854 5256
rect -29907 5220 -29610 5238
rect -29592 5220 -29313 5238
rect -29907 5193 -29880 5220
rect -30357 5175 -29880 5193
rect -30357 5121 -30339 5175
rect -30204 5121 -30186 5175
rect -29907 5166 -29880 5175
rect -29331 5184 -29313 5220
rect -29178 5184 -29160 5238
rect -28881 5229 -28854 5238
rect -30303 5040 -30285 5094
rect -30141 5040 -30123 5103
rect -29979 5049 -29889 5076
rect -29979 5040 -29961 5049
rect -30303 5022 -29961 5040
rect -29835 5040 -29808 5130
rect -29277 5103 -29259 5157
rect -29115 5103 -29097 5166
rect -28953 5112 -28863 5139
rect -28953 5103 -28935 5112
rect -29277 5085 -28935 5103
rect -28809 5103 -28782 5193
rect -29115 5049 -29097 5085
rect -30141 4986 -30123 5022
rect -28881 5040 -28854 5067
rect -29907 4977 -29880 5004
rect -29331 5004 -29313 5022
rect -28881 5022 -28782 5040
rect -28881 5004 -28845 5022
rect -29331 4986 -28989 5004
rect -28971 4986 -28845 5004
rect -29331 4977 -29313 4986
rect -30357 4941 -30339 4959
rect -29907 4959 -29529 4977
rect -29511 4959 -29313 4977
rect -29907 4941 -29871 4959
rect -31104 4923 -29871 4941
rect -31104 3006 -31086 4923
rect -29889 4590 -29871 4923
rect -29691 4797 -29610 4815
rect -29592 4797 -29421 4815
rect -29691 4761 -29673 4797
rect -29466 4761 -29448 4797
rect -29538 4680 -29520 4734
rect -29412 4680 -29394 4734
rect -29628 4662 -29439 4680
rect -29412 4662 -29403 4680
rect -29628 4635 -29610 4662
rect -29538 4635 -29520 4662
rect -29412 4635 -29394 4662
rect -29682 4590 -29664 4617
rect -29592 4590 -29574 4617
rect -29466 4590 -29448 4617
rect -29889 4572 -29448 4590
rect -29574 4365 -29538 4383
rect -30438 4149 -30222 4185
rect -30186 4149 -30006 4185
rect -29628 4149 -29412 4185
rect -29376 4149 -29196 4185
rect -28746 4149 -28530 4185
rect -28494 4149 -28314 4185
rect -30438 4077 -30222 4113
rect -30186 4077 -30051 4113
rect -30087 4041 -30051 4077
rect -30600 3978 -30474 4014
rect -30438 3978 -30222 4014
rect -30600 3879 -30564 3978
rect -30087 3942 -30051 4023
rect -30438 3906 -30222 3942
rect -30186 3906 -30051 3942
rect -30042 3879 -30006 4149
rect -29628 4077 -29412 4113
rect -29376 4077 -29241 4113
rect -29277 4041 -29241 4077
rect -30600 3843 -30375 3879
rect -30780 3807 -30726 3825
rect -30600 3789 -30474 3825
rect -30726 3753 -30708 3762
rect -30726 3744 -30699 3753
rect -30600 3726 -30564 3753
rect -30411 3744 -30375 3843
rect -30357 3843 -30006 3879
rect -29790 3978 -29664 4014
rect -29628 3978 -29412 4014
rect -29790 3879 -29754 3978
rect -29277 3942 -29241 4023
rect -29628 3906 -29412 3942
rect -29376 3906 -29241 3942
rect -29232 3879 -29196 4149
rect -28746 4077 -28530 4113
rect -28494 4077 -28359 4113
rect -28395 4050 -28359 4077
rect -29790 3843 -29565 3879
rect -30357 3834 -30321 3843
rect -30186 3789 -30069 3825
rect -30537 3735 -30528 3744
rect -30555 3726 -30528 3735
rect -30753 3708 -30564 3726
rect -30438 3708 -30222 3744
rect -30105 3726 -30069 3753
rect -29790 3789 -29664 3825
rect -30105 3708 -29979 3726
rect -29952 3717 -29898 3735
rect -30753 3006 -30735 3708
rect -30600 3699 -30564 3708
rect -30105 3699 -30069 3708
rect -30600 3627 -30474 3663
rect -30186 3627 -30069 3663
rect -30438 3546 -30222 3582
rect -30357 3519 -30321 3546
rect -29997 3258 -29979 3708
rect -29790 3699 -29754 3753
rect -29601 3744 -29565 3843
rect -29547 3843 -29196 3879
rect -28908 3978 -28782 4014
rect -28746 3978 -28530 4014
rect -28908 3879 -28872 3978
rect -28395 3942 -28359 4005
rect -28746 3906 -28530 3942
rect -28494 3906 -28359 3942
rect -28350 3879 -28314 4149
rect -28908 3843 -28683 3879
rect -29547 3834 -29511 3843
rect -29376 3789 -29259 3825
rect -29628 3708 -29412 3744
rect -29295 3735 -29259 3753
rect -28908 3789 -28782 3825
rect -28908 3735 -28872 3753
rect -28719 3744 -28683 3843
rect -28665 3843 -28314 3879
rect -28665 3834 -28629 3843
rect -28494 3789 -28377 3825
rect -29295 3717 -29178 3735
rect -29718 3699 -29700 3708
rect -29295 3699 -29259 3717
rect -29790 3627 -29664 3663
rect -29718 3348 -29700 3627
rect -29376 3627 -29259 3663
rect -29628 3546 -29412 3582
rect -29547 3519 -29511 3546
rect -29718 3330 -29538 3348
rect -29196 3321 -29178 3717
rect -29070 3708 -29043 3735
rect -28917 3717 -28872 3735
rect -28908 3699 -28872 3717
rect -28746 3708 -28530 3744
rect -28413 3735 -28377 3753
rect -28413 3717 -28368 3735
rect -28836 3699 -28809 3708
rect -28413 3699 -28377 3717
rect -28908 3627 -28782 3663
rect -28494 3627 -28377 3663
rect -28881 3420 -28863 3627
rect -28746 3546 -28530 3582
rect -28665 3519 -28629 3546
rect -28971 3402 -28863 3420
rect -28350 3411 -28332 3717
rect -28881 3348 -28350 3366
rect -28881 3321 -28854 3348
rect -29331 3303 -28854 3321
rect -29907 3285 -29610 3303
rect -29592 3285 -29313 3303
rect -29907 3258 -29880 3285
rect -30357 3240 -29880 3258
rect -30357 3186 -30339 3240
rect -30204 3186 -30186 3240
rect -29907 3231 -29880 3240
rect -29331 3249 -29313 3285
rect -29178 3249 -29160 3303
rect -28881 3294 -28854 3303
rect -30303 3105 -30285 3159
rect -30141 3105 -30123 3168
rect -29979 3114 -29889 3141
rect -29979 3105 -29961 3114
rect -30303 3087 -29961 3105
rect -29835 3105 -29808 3195
rect -29277 3168 -29259 3222
rect -29115 3168 -29097 3231
rect -28953 3177 -28863 3204
rect -28953 3168 -28935 3177
rect -29277 3150 -28935 3168
rect -28809 3168 -28782 3258
rect -29115 3114 -29097 3150
rect -30141 3051 -30123 3087
rect -28881 3105 -28854 3132
rect -29907 3042 -29880 3069
rect -29331 3069 -29313 3087
rect -28881 3087 -28782 3105
rect -28881 3069 -28845 3087
rect -29331 3051 -28989 3069
rect -28971 3051 -28845 3069
rect -29331 3042 -29313 3051
rect -30357 3006 -30339 3024
rect -29907 3024 -29529 3042
rect -29511 3024 -29313 3042
rect -29907 3006 -29871 3024
rect -31104 2988 -29871 3006
rect -29889 2655 -29871 2988
rect -29691 2862 -29610 2880
rect -29592 2862 -29421 2880
rect -29691 2826 -29673 2862
rect -29466 2826 -29448 2862
rect -29538 2745 -29520 2799
rect -29412 2745 -29394 2799
rect -27990 2745 -27972 5436
rect -29628 2727 -29439 2745
rect -29412 2727 -27972 2745
rect -29628 2700 -29610 2727
rect -29538 2700 -29520 2727
rect -29412 2700 -29394 2727
rect -29682 2655 -29664 2682
rect -29592 2655 -29574 2682
rect -29466 2655 -29448 2682
rect -30402 2637 -29448 2655
rect -37332 2340 -33507 2349
rect -30402 2340 -30384 2637
rect -37332 2322 -30384 2340
rect -37332 -13428 -37296 2322
rect -36801 -1341 -36783 1035
rect -30402 45 -30384 2322
rect -30078 459 -29862 495
rect -29826 459 -29646 495
rect -30078 387 -29862 423
rect -29826 387 -29691 423
rect -30240 288 -30114 324
rect -30078 288 -29862 324
rect -29727 306 -29691 387
rect -30240 189 -30204 288
rect -29727 270 -29718 306
rect -29727 252 -29691 270
rect -30078 216 -29862 252
rect -29826 216 -29691 252
rect -29682 189 -29646 459
rect -30240 153 -30015 189
rect -30240 99 -30114 135
rect -30240 45 -30204 63
rect -30051 54 -30015 153
rect -29997 153 -29646 189
rect -29610 450 -29322 468
rect -29997 144 -29961 153
rect -29826 99 -29709 135
rect -30402 27 -30204 45
rect -30825 -99 -30744 -81
rect -33435 -234 -33201 -216
rect -33435 -261 -33408 -234
rect -34236 -279 -33408 -261
rect -34236 -1026 -34218 -279
rect -33885 -333 -33867 -279
rect -33732 -333 -33714 -279
rect -33435 -288 -33408 -279
rect -33831 -414 -33813 -360
rect -33669 -414 -33651 -351
rect -33363 -369 -33336 -324
rect -33507 -405 -33417 -378
rect -33363 -396 -33354 -369
rect -33507 -414 -33489 -405
rect -33831 -432 -33489 -414
rect -33363 -414 -33336 -396
rect -33669 -468 -33651 -432
rect -33435 -477 -33408 -450
rect -33885 -513 -33867 -495
rect -33435 -495 -33336 -477
rect -33435 -513 -33399 -495
rect -33993 -531 -33399 -513
rect -33993 -1008 -33975 -531
rect -33696 -594 -33678 -585
rect -33219 -711 -33201 -234
rect -30402 -261 -30384 27
rect -30240 9 -30204 27
rect -30078 18 -29862 54
rect -29745 45 -29709 63
rect -29610 45 -29583 450
rect -29520 441 -29484 450
rect -29511 396 -29484 441
rect -29439 315 -29412 360
rect -29439 288 -29376 315
rect -29439 270 -29412 288
rect -29511 207 -29484 234
rect -29745 18 -29583 45
rect -29538 189 -29448 207
rect -29745 9 -29709 18
rect -29970 -27 -29943 -9
rect -30240 -63 -30114 -27
rect -29826 -63 -29709 -27
rect -30339 -99 -30285 -81
rect -30078 -144 -29862 -108
rect -29997 -171 -29961 -144
rect -29538 -261 -29520 189
rect -30402 -279 -29520 -261
rect -29340 153 -29322 450
rect -28305 180 -28206 189
rect -28305 153 -28278 180
rect -29340 135 -28431 153
rect -28404 135 -28278 153
rect -30618 -351 -30465 -333
rect -33435 -729 -33201 -711
rect -33435 -756 -33408 -729
rect -33885 -774 -33408 -756
rect -33885 -828 -33867 -774
rect -33732 -828 -33714 -774
rect -33435 -783 -33408 -774
rect -33831 -909 -33813 -855
rect -33669 -909 -33651 -846
rect -33363 -864 -33336 -819
rect -33507 -900 -33417 -873
rect -33363 -891 -33354 -864
rect -33507 -909 -33489 -900
rect -33831 -927 -33489 -909
rect -33363 -909 -33336 -891
rect -33669 -963 -33651 -927
rect -33435 -972 -33408 -945
rect -33885 -1008 -33867 -990
rect -33435 -990 -33336 -972
rect -33435 -1008 -33399 -990
rect -33993 -1026 -33399 -1008
rect -34461 -1044 -34191 -1026
rect -34461 -1080 -34443 -1044
rect -34236 -1080 -34218 -1044
rect -34308 -1161 -34290 -1107
rect -34398 -1179 -34209 -1161
rect -34398 -1206 -34380 -1179
rect -34308 -1206 -34290 -1179
rect -34182 -1206 -34164 -1107
rect -34452 -1251 -34434 -1224
rect -34362 -1251 -34344 -1224
rect -34236 -1251 -34218 -1224
rect -33993 -1251 -33975 -1026
rect -33219 -1125 -33201 -729
rect -33435 -1143 -33201 -1125
rect -33435 -1170 -33408 -1143
rect -34470 -1269 -33975 -1251
rect -33885 -1188 -33408 -1170
rect -33885 -1242 -33867 -1188
rect -33732 -1242 -33714 -1188
rect -33435 -1197 -33408 -1188
rect -33993 -1422 -33975 -1269
rect -33831 -1323 -33813 -1269
rect -33669 -1323 -33651 -1260
rect -33363 -1278 -33336 -1233
rect -33507 -1314 -33417 -1287
rect -33363 -1305 -33354 -1278
rect -33507 -1323 -33489 -1314
rect -33831 -1341 -33489 -1323
rect -33363 -1323 -33336 -1305
rect -33669 -1377 -33651 -1341
rect -33435 -1386 -33408 -1359
rect -33885 -1422 -33867 -1404
rect -33435 -1404 -33336 -1386
rect -33435 -1422 -33399 -1404
rect -33993 -1440 -33399 -1422
rect -35361 -1557 -35352 -1539
rect -33993 -1953 -33975 -1440
rect -33696 -1530 -33678 -1494
rect -33219 -1656 -33201 -1143
rect -33435 -1674 -33201 -1656
rect -33435 -1701 -33408 -1674
rect -33885 -1719 -33408 -1701
rect -33885 -1773 -33867 -1719
rect -33732 -1773 -33714 -1719
rect -33435 -1728 -33408 -1719
rect -33831 -1854 -33813 -1800
rect -33669 -1854 -33651 -1791
rect -33363 -1809 -33336 -1764
rect -33507 -1845 -33417 -1818
rect -33363 -1836 -33354 -1809
rect -33507 -1854 -33489 -1845
rect -33831 -1872 -33489 -1854
rect -33363 -1854 -33336 -1836
rect -33669 -1908 -33651 -1872
rect -33435 -1917 -33408 -1890
rect -33885 -1953 -33867 -1935
rect -33435 -1935 -33336 -1917
rect -33435 -1953 -33399 -1935
rect -33993 -1971 -33399 -1953
rect -35262 -2106 -35235 -2088
rect -33993 -2520 -33975 -1971
rect -33696 -2079 -33678 -2052
rect -33219 -2223 -33201 -1674
rect -33435 -2241 -33201 -2223
rect -33435 -2268 -33408 -2241
rect -33930 -2286 -33408 -2268
rect -33885 -2340 -33867 -2286
rect -33732 -2340 -33714 -2286
rect -33435 -2295 -33408 -2286
rect -33831 -2421 -33813 -2367
rect -33669 -2421 -33651 -2358
rect -33363 -2376 -33336 -2331
rect -33507 -2412 -33417 -2385
rect -33363 -2403 -33354 -2376
rect -33507 -2421 -33489 -2412
rect -33831 -2439 -33489 -2421
rect -33363 -2421 -33336 -2403
rect -33669 -2475 -33651 -2439
rect -33435 -2484 -33408 -2457
rect -33885 -2520 -33867 -2502
rect -33435 -2502 -33336 -2484
rect -33435 -2520 -33399 -2502
rect -33993 -2538 -33399 -2520
rect -34605 -2655 -34596 -2628
rect -33993 -3015 -33975 -2538
rect -33696 -2628 -33678 -2601
rect -33219 -2718 -33201 -2241
rect -33435 -2736 -33201 -2718
rect -33435 -2763 -33408 -2736
rect -33885 -2781 -33408 -2763
rect -33885 -2835 -33867 -2781
rect -33732 -2835 -33714 -2781
rect -33435 -2790 -33408 -2781
rect -33831 -2916 -33813 -2862
rect -33669 -2916 -33651 -2853
rect -33363 -2871 -33336 -2826
rect -33507 -2907 -33417 -2880
rect -33363 -2898 -33345 -2871
rect -33507 -2916 -33489 -2907
rect -33831 -2934 -33489 -2916
rect -33363 -2916 -33336 -2898
rect -33669 -2970 -33651 -2934
rect -33435 -2979 -33408 -2952
rect -33885 -3015 -33867 -2997
rect -33435 -2997 -33336 -2979
rect -33435 -3015 -33399 -2997
rect -33993 -3033 -33399 -3015
rect -34776 -3123 -34758 -3087
rect -33993 -3258 -33975 -3033
rect -33696 -3087 -33678 -3078
rect -33219 -3132 -33201 -2736
rect -33435 -3150 -33201 -3132
rect -33435 -3177 -33408 -3150
rect -34029 -3276 -33975 -3258
rect -33885 -3195 -33408 -3177
rect -33885 -3249 -33867 -3195
rect -33732 -3249 -33714 -3195
rect -33435 -3204 -33408 -3195
rect -33993 -3429 -33975 -3276
rect -33831 -3330 -33813 -3276
rect -33669 -3330 -33651 -3267
rect -33363 -3285 -33336 -3240
rect -33507 -3321 -33417 -3294
rect -33363 -3312 -33345 -3285
rect -33507 -3330 -33489 -3321
rect -33831 -3348 -33489 -3330
rect -33363 -3330 -33336 -3312
rect -33669 -3384 -33651 -3348
rect -33435 -3393 -33408 -3366
rect -33885 -3429 -33867 -3411
rect -33435 -3411 -33336 -3393
rect -33435 -3429 -33399 -3411
rect -33993 -3447 -33399 -3429
rect -34956 -3627 -34947 -3600
rect -33993 -3960 -33975 -3447
rect -33696 -3537 -33678 -3519
rect -33219 -3663 -33201 -3150
rect -31365 -882 -30717 -864
rect -33435 -3681 -33174 -3663
rect -33435 -3708 -33408 -3681
rect -33885 -3726 -33408 -3708
rect -33885 -3780 -33867 -3726
rect -33732 -3780 -33714 -3726
rect -33435 -3735 -33408 -3726
rect -33831 -3861 -33813 -3807
rect -33669 -3861 -33651 -3798
rect -33363 -3816 -33336 -3771
rect -33507 -3852 -33417 -3825
rect -33363 -3843 -33345 -3816
rect -33507 -3861 -33489 -3852
rect -33831 -3879 -33489 -3861
rect -33363 -3861 -33336 -3843
rect -33669 -3915 -33651 -3879
rect -33435 -3924 -33408 -3897
rect -33885 -3960 -33867 -3942
rect -33435 -3942 -33336 -3924
rect -33435 -3960 -33399 -3942
rect -33993 -3978 -33399 -3960
rect -35127 -4131 -35064 -4104
rect -33993 -8100 -33975 -3978
rect -33696 -4050 -33678 -4041
rect -33201 -8073 -33174 -3681
rect -31716 -3843 -31698 -3816
rect -31797 -3852 -31698 -3843
rect -31680 -3852 -31644 -3816
rect -31365 -5670 -31338 -882
rect -30402 -900 -30384 -279
rect -30078 -486 -29862 -450
rect -29826 -486 -29646 -450
rect -29340 -477 -29322 135
rect -29142 90 -29115 135
rect -28755 81 -28737 135
rect -28602 81 -28584 135
rect -28305 126 -28278 135
rect -29070 -36 -29043 54
rect -28701 0 -28683 54
rect -28539 0 -28521 63
rect -28233 45 -28206 90
rect -28377 9 -28287 36
rect -28233 18 -27045 45
rect -28377 0 -28359 9
rect -28701 -18 -28359 0
rect -28233 0 -28206 18
rect -28539 -54 -28521 -18
rect -29142 -99 -29115 -72
rect -28305 -63 -28278 -36
rect -28755 -99 -28737 -81
rect -28305 -81 -28206 -63
rect -28305 -99 -28269 -81
rect -29124 -117 -28269 -99
rect -30078 -558 -29862 -522
rect -29826 -558 -29691 -522
rect -30240 -657 -30114 -621
rect -30078 -657 -29862 -621
rect -29727 -639 -29691 -558
rect -30240 -756 -30204 -657
rect -29727 -675 -29718 -639
rect -29727 -693 -29691 -675
rect -30078 -729 -29862 -693
rect -29826 -729 -29691 -693
rect -29682 -756 -29646 -486
rect -30240 -792 -30015 -756
rect -30240 -846 -30114 -810
rect -30240 -900 -30204 -882
rect -30051 -891 -30015 -792
rect -29997 -792 -29646 -756
rect -29610 -495 -29322 -477
rect -29997 -801 -29961 -792
rect -29826 -846 -29709 -810
rect -30402 -918 -30204 -900
rect -30942 -1044 -30915 -1026
rect -30402 -1206 -30384 -918
rect -30240 -936 -30204 -918
rect -30078 -927 -29862 -891
rect -29745 -900 -29709 -882
rect -29610 -900 -29583 -495
rect -29520 -504 -29484 -495
rect -29511 -549 -29484 -504
rect -29439 -630 -29412 -585
rect -29439 -657 -29385 -630
rect -29340 -657 -29322 -495
rect -27882 -522 -27864 -432
rect -28377 -630 -28278 -621
rect -27549 -630 -27108 -612
rect -28377 -657 -28350 -630
rect -27549 -657 -27522 -630
rect -29439 -675 -29412 -657
rect -29340 -675 -27522 -657
rect -29511 -738 -29484 -711
rect -29745 -927 -29583 -900
rect -29538 -756 -29475 -738
rect -29457 -756 -29421 -738
rect -29745 -936 -29709 -927
rect -29970 -972 -29943 -954
rect -30240 -1008 -30114 -972
rect -29826 -1008 -29709 -972
rect -30339 -1044 -30285 -1026
rect -30078 -1089 -29862 -1053
rect -29997 -1116 -29961 -1089
rect -29538 -1206 -29520 -756
rect -30402 -1224 -29520 -1206
rect -30402 -1917 -30384 -1224
rect -29340 -1431 -29322 -675
rect -29160 -720 -29133 -675
rect -28827 -729 -28809 -675
rect -28674 -729 -28656 -675
rect -28377 -684 -28350 -675
rect -29088 -846 -29061 -756
rect -28773 -810 -28755 -756
rect -28611 -810 -28593 -747
rect -28449 -801 -28359 -774
rect -28449 -810 -28431 -801
rect -28773 -828 -28431 -810
rect -28305 -810 -28278 -720
rect -27999 -729 -27981 -675
rect -27846 -729 -27828 -675
rect -27549 -684 -27522 -675
rect -27126 -684 -27108 -630
rect -28611 -864 -28593 -828
rect -29160 -909 -29133 -882
rect -27945 -810 -27927 -756
rect -27783 -810 -27765 -747
rect -27477 -765 -27450 -720
rect -27126 -702 -26676 -684
rect -27126 -738 -27108 -702
rect -26721 -738 -26703 -702
rect -27621 -801 -27531 -774
rect -27477 -792 -27270 -765
rect -27621 -810 -27603 -801
rect -27945 -828 -27603 -810
rect -27477 -810 -27450 -792
rect -28377 -873 -28350 -846
rect -27783 -864 -27765 -828
rect -28827 -909 -28809 -891
rect -28377 -891 -28278 -873
rect -27288 -801 -27270 -792
rect -27288 -819 -27090 -801
rect -26793 -819 -26775 -765
rect -26667 -819 -26649 -765
rect -27063 -837 -26694 -819
rect -26667 -837 -26622 -819
rect -27549 -873 -27522 -846
rect -27063 -864 -27045 -837
rect -26973 -864 -26955 -837
rect -26883 -864 -26865 -837
rect -26793 -864 -26775 -837
rect -26667 -864 -26649 -837
rect -28377 -909 -28341 -891
rect -27999 -909 -27981 -891
rect -27549 -891 -27450 -873
rect -27549 -909 -27513 -891
rect -27126 -909 -27108 -882
rect -27027 -909 -27009 -882
rect -26937 -909 -26919 -882
rect -26847 -909 -26829 -882
rect -26721 -909 -26703 -882
rect -29124 -927 -26703 -909
rect -29340 -1458 -27846 -1431
rect -30078 -1503 -29862 -1467
rect -29826 -1503 -29646 -1467
rect -29340 -1494 -29322 -1458
rect -30078 -1575 -29862 -1539
rect -29826 -1575 -29691 -1539
rect -30240 -1674 -30114 -1638
rect -30078 -1674 -29862 -1638
rect -29727 -1656 -29691 -1575
rect -30240 -1773 -30204 -1674
rect -29727 -1692 -29718 -1656
rect -29727 -1710 -29691 -1692
rect -30078 -1746 -29862 -1710
rect -29826 -1746 -29691 -1710
rect -29682 -1773 -29646 -1503
rect -30240 -1809 -30015 -1773
rect -30240 -1863 -30114 -1827
rect -30240 -1917 -30204 -1899
rect -30051 -1908 -30015 -1809
rect -29997 -1809 -29646 -1773
rect -29610 -1503 -29322 -1494
rect -28674 -1503 -28647 -1458
rect -29610 -1512 -29079 -1503
rect -29997 -1818 -29961 -1809
rect -29826 -1863 -29709 -1827
rect -30402 -1935 -30204 -1917
rect -31077 -2061 -30924 -2043
rect -31365 -5688 -31131 -5670
rect -31284 -6687 -31266 -6606
rect -31419 -6813 -31311 -6786
rect -33417 -8091 -33174 -8073
rect -33993 -8127 -33957 -8100
rect -33417 -8118 -33390 -8091
rect -35676 -8451 -35658 -8424
rect -33975 -8370 -33957 -8127
rect -33867 -8136 -33390 -8118
rect -33201 -8127 -33174 -8091
rect -33867 -8190 -33849 -8136
rect -33714 -8190 -33696 -8136
rect -33417 -8145 -33390 -8136
rect -33813 -8271 -33795 -8217
rect -33651 -8271 -33633 -8208
rect -33345 -8226 -33318 -8181
rect -33489 -8262 -33399 -8235
rect -33345 -8253 -33336 -8226
rect -33489 -8271 -33471 -8262
rect -33813 -8289 -33471 -8271
rect -33345 -8271 -33318 -8253
rect -33651 -8325 -33633 -8289
rect -33417 -8334 -33390 -8307
rect -33867 -8370 -33849 -8352
rect -33417 -8352 -33318 -8334
rect -33417 -8370 -33381 -8352
rect -33975 -8388 -33381 -8370
rect -34173 -8478 -34164 -8460
rect -33975 -8865 -33957 -8388
rect -33678 -8451 -33660 -8433
rect -33192 -8568 -33174 -8127
rect -33417 -8586 -33174 -8568
rect -33417 -8613 -33390 -8586
rect -33867 -8631 -33390 -8613
rect -33867 -8685 -33849 -8631
rect -33714 -8685 -33696 -8631
rect -33417 -8640 -33390 -8631
rect -33813 -8766 -33795 -8712
rect -33651 -8766 -33633 -8703
rect -33345 -8721 -33318 -8676
rect -33489 -8757 -33399 -8730
rect -33345 -8748 -33327 -8721
rect -33489 -8766 -33471 -8757
rect -33813 -8784 -33471 -8766
rect -33345 -8766 -33318 -8748
rect -33651 -8820 -33633 -8784
rect -33417 -8829 -33390 -8802
rect -33867 -8865 -33849 -8847
rect -33417 -8847 -33318 -8829
rect -33417 -8865 -33381 -8847
rect -33975 -8883 -33381 -8865
rect -35523 -8928 -35505 -8919
rect -34236 -8973 -34218 -8964
rect -33975 -9279 -33957 -8883
rect -33192 -8982 -33174 -8586
rect -31230 -8721 -31212 -5688
rect -31077 -6606 -31050 -2061
rect -30402 -2223 -30384 -1935
rect -30240 -1953 -30204 -1935
rect -30078 -1944 -29862 -1908
rect -29745 -1917 -29709 -1899
rect -29610 -1917 -29583 -1512
rect -29520 -1521 -29484 -1512
rect -29511 -1566 -29484 -1521
rect -29340 -1521 -29151 -1512
rect -29439 -1692 -29412 -1602
rect -29511 -1755 -29484 -1728
rect -29745 -1944 -29583 -1917
rect -29538 -1773 -29457 -1755
rect -29745 -1953 -29709 -1944
rect -30240 -2025 -30114 -1989
rect -29943 -1998 -29925 -1980
rect -29826 -2025 -29709 -1989
rect -30339 -2061 -30285 -2043
rect -30078 -2106 -29862 -2070
rect -29997 -2133 -29961 -2106
rect -29916 -2169 -29898 -2151
rect -29538 -2223 -29520 -1773
rect -30402 -2241 -29520 -2223
rect -30789 -2340 -30771 -2322
rect -30708 -2403 -30483 -2385
rect -30402 -3213 -30384 -2241
rect -29340 -2727 -29322 -1521
rect -29178 -1566 -29151 -1521
rect -28548 -1503 -28521 -1458
rect -28404 -1503 -28377 -1458
rect -28611 -1584 -28584 -1539
rect -28278 -1503 -28251 -1458
rect -28485 -1584 -28458 -1539
rect -28152 -1503 -28125 -1458
rect -28341 -1584 -28314 -1539
rect -27882 -1494 -27855 -1458
rect -28215 -1584 -28188 -1539
rect -28080 -1584 -28053 -1539
rect -27819 -1584 -27792 -1539
rect -26946 -1584 -26928 -1233
rect -29106 -1647 -29079 -1602
rect -28881 -1629 -28656 -1602
rect -28611 -1611 -27855 -1584
rect -27819 -1611 -26928 -1584
rect -28881 -1647 -28863 -1629
rect -28278 -1647 -28251 -1620
rect -29106 -1674 -28863 -1647
rect -28053 -1674 -28026 -1611
rect -27819 -1674 -27792 -1611
rect -29106 -1692 -29079 -1674
rect -29178 -1755 -29151 -1728
rect -28674 -1746 -28647 -1701
rect -27882 -1746 -27855 -1701
rect -28674 -1755 -27855 -1746
rect -29187 -1773 -29178 -1755
rect -29142 -1773 -27855 -1755
rect -29340 -2754 -27999 -2727
rect -30078 -2799 -29862 -2763
rect -29826 -2799 -29646 -2763
rect -29340 -2790 -29322 -2754
rect -30078 -2871 -29862 -2835
rect -29826 -2871 -29691 -2835
rect -30240 -2970 -30114 -2934
rect -30078 -2970 -29862 -2934
rect -29727 -2952 -29691 -2871
rect -30240 -3069 -30204 -2970
rect -29727 -2988 -29718 -2952
rect -29727 -3006 -29691 -2988
rect -30078 -3042 -29862 -3006
rect -29826 -3042 -29691 -3006
rect -29682 -3069 -29646 -2799
rect -30240 -3105 -30015 -3069
rect -30240 -3159 -30114 -3123
rect -30240 -3213 -30204 -3195
rect -30051 -3204 -30015 -3105
rect -29997 -3105 -29646 -3069
rect -29610 -2808 -29133 -2790
rect -28827 -2799 -28800 -2754
rect -29997 -3114 -29961 -3105
rect -29826 -3159 -29709 -3123
rect -30402 -3231 -30204 -3213
rect -30402 -3519 -30384 -3231
rect -30240 -3249 -30204 -3231
rect -30078 -3240 -29862 -3204
rect -29745 -3213 -29709 -3195
rect -29610 -3195 -29583 -2808
rect -29520 -2817 -29484 -2808
rect -29241 -2817 -29205 -2808
rect -29511 -2862 -29484 -2817
rect -29232 -2862 -29205 -2817
rect -28701 -2799 -28674 -2754
rect -28557 -2799 -28530 -2754
rect -29439 -2943 -29412 -2898
rect -28764 -2880 -28737 -2835
rect -28431 -2799 -28404 -2754
rect -28638 -2880 -28611 -2835
rect -28305 -2799 -28278 -2754
rect -28494 -2880 -28467 -2835
rect -28035 -2790 -28008 -2754
rect -28368 -2880 -28341 -2835
rect -28233 -2880 -28206 -2835
rect -27972 -2880 -27945 -2835
rect -26856 -2880 -26838 -1647
rect -29160 -2943 -29133 -2898
rect -28971 -2925 -28809 -2898
rect -28764 -2907 -28008 -2880
rect -27972 -2907 -26838 -2880
rect -28971 -2943 -28953 -2925
rect -29439 -2970 -29385 -2943
rect -29439 -2988 -29412 -2970
rect -29160 -2970 -28953 -2943
rect -28206 -2970 -28179 -2907
rect -27972 -2970 -27945 -2907
rect -29160 -2988 -29133 -2970
rect -29511 -3051 -29484 -3024
rect -29232 -3051 -29205 -3024
rect -28827 -3042 -28800 -2997
rect -28035 -3042 -28008 -2997
rect -28827 -3051 -28008 -3042
rect -29745 -3240 -29610 -3213
rect -29538 -3069 -28008 -3051
rect -29745 -3249 -29709 -3240
rect -29943 -3285 -29925 -3276
rect -30240 -3321 -30114 -3285
rect -29826 -3321 -29709 -3285
rect -30078 -3402 -29862 -3366
rect -29997 -3429 -29961 -3402
rect -29538 -3519 -29520 -3069
rect -30402 -3537 -29520 -3519
rect -30789 -3663 -30762 -3645
rect -30987 -3744 -30798 -3726
rect -30402 -4284 -30384 -3537
rect -29790 -3636 -29772 -3627
rect -30078 -3870 -29862 -3834
rect -29826 -3870 -29646 -3834
rect -30078 -3942 -29862 -3906
rect -29826 -3942 -29691 -3906
rect -30240 -4041 -30114 -4005
rect -30078 -4041 -29862 -4005
rect -29727 -4023 -29691 -3942
rect -30240 -4140 -30204 -4041
rect -29727 -4059 -29718 -4023
rect -29727 -4077 -29691 -4059
rect -30078 -4113 -29862 -4077
rect -29826 -4113 -29691 -4077
rect -29682 -4140 -29646 -3870
rect -30240 -4176 -30015 -4140
rect -30240 -4230 -30114 -4194
rect -30240 -4284 -30204 -4266
rect -30051 -4275 -30015 -4176
rect -29997 -4176 -29646 -4140
rect -29583 -3879 -29322 -3861
rect -29520 -3888 -29484 -3879
rect -29997 -4185 -29961 -4176
rect -29826 -4230 -29709 -4194
rect -30402 -4302 -30204 -4284
rect -30402 -4590 -30384 -4302
rect -30240 -4320 -30204 -4302
rect -30078 -4311 -29862 -4275
rect -29745 -4284 -29709 -4266
rect -29610 -4284 -29583 -3915
rect -29511 -3933 -29484 -3888
rect -29439 -4014 -29412 -3969
rect -29439 -4041 -29376 -4014
rect -29439 -4059 -29412 -4041
rect -29511 -4122 -29484 -4095
rect -29745 -4311 -29583 -4284
rect -29538 -4140 -29448 -4122
rect -29745 -4320 -29709 -4311
rect -29970 -4356 -29943 -4338
rect -30240 -4392 -30114 -4356
rect -29826 -4392 -29709 -4356
rect -30078 -4473 -29862 -4437
rect -29997 -4500 -29961 -4473
rect -29538 -4590 -29520 -4140
rect -30402 -4608 -29520 -4590
rect -29340 -4176 -29322 -3879
rect -28305 -4149 -28206 -4140
rect -28305 -4176 -28278 -4149
rect -29340 -4194 -28278 -4176
rect -30879 -4680 -30852 -4662
rect -30402 -5229 -30384 -4608
rect -30078 -4815 -29862 -4779
rect -29826 -4815 -29646 -4779
rect -29340 -4806 -29322 -4194
rect -29142 -4239 -29115 -4194
rect -28755 -4248 -28737 -4194
rect -28602 -4248 -28584 -4194
rect -28305 -4203 -28278 -4194
rect -29070 -4365 -29043 -4275
rect -28701 -4329 -28683 -4275
rect -28539 -4329 -28521 -4266
rect -28233 -4284 -28206 -4239
rect -28377 -4320 -28287 -4293
rect -28233 -4311 -27045 -4284
rect -28377 -4329 -28359 -4320
rect -28701 -4347 -28359 -4329
rect -28233 -4329 -28206 -4311
rect -28539 -4383 -28521 -4347
rect -29142 -4428 -29115 -4401
rect -28305 -4392 -28278 -4365
rect -28755 -4428 -28737 -4410
rect -28305 -4410 -28206 -4392
rect -28305 -4428 -28269 -4410
rect -29124 -4446 -28269 -4428
rect -30078 -4887 -29862 -4851
rect -29826 -4887 -29691 -4851
rect -30240 -4986 -30114 -4950
rect -30078 -4986 -29862 -4950
rect -29727 -4968 -29691 -4887
rect -30240 -5085 -30204 -4986
rect -29727 -5004 -29718 -4968
rect -29727 -5022 -29691 -5004
rect -30078 -5058 -29862 -5022
rect -29826 -5058 -29691 -5022
rect -29682 -5085 -29646 -4815
rect -30240 -5121 -30015 -5085
rect -30240 -5175 -30114 -5139
rect -30240 -5229 -30204 -5211
rect -30051 -5220 -30015 -5121
rect -29997 -5121 -29646 -5085
rect -29610 -4824 -29322 -4806
rect -29997 -5130 -29961 -5121
rect -29826 -5175 -29709 -5139
rect -30402 -5247 -30204 -5229
rect -30960 -5616 -30942 -5409
rect -30402 -5535 -30384 -5247
rect -30240 -5265 -30204 -5247
rect -30078 -5256 -29862 -5220
rect -29745 -5229 -29709 -5211
rect -29610 -5229 -29583 -4824
rect -29520 -4833 -29484 -4824
rect -29511 -4878 -29484 -4833
rect -29439 -4959 -29412 -4914
rect -29439 -4986 -29385 -4959
rect -29340 -4986 -29322 -4824
rect -27882 -4851 -27864 -4761
rect -28377 -4959 -28278 -4950
rect -27549 -4959 -27108 -4941
rect -28377 -4986 -28350 -4959
rect -27549 -4986 -27522 -4959
rect -29439 -5004 -29412 -4986
rect -29340 -5004 -27522 -4986
rect -29511 -5067 -29484 -5040
rect -29745 -5256 -29583 -5229
rect -29538 -5085 -29475 -5067
rect -29457 -5085 -29421 -5067
rect -29745 -5265 -29709 -5256
rect -29970 -5301 -29943 -5283
rect -30240 -5337 -30114 -5301
rect -29826 -5337 -29709 -5301
rect -30240 -5508 -30213 -5373
rect -30078 -5418 -29862 -5382
rect -29997 -5445 -29961 -5418
rect -29538 -5535 -29520 -5085
rect -31167 -7965 -31149 -7947
rect -31500 -8748 -31212 -8721
rect -33417 -9000 -33174 -8982
rect -33417 -9027 -33390 -9000
rect -33867 -9045 -33390 -9027
rect -33867 -9099 -33849 -9045
rect -33714 -9099 -33696 -9045
rect -33417 -9054 -33390 -9045
rect -33813 -9180 -33795 -9126
rect -33651 -9180 -33633 -9117
rect -33489 -9171 -33399 -9144
rect -33489 -9180 -33471 -9171
rect -33813 -9198 -33471 -9180
rect -33345 -9180 -33318 -9090
rect -33651 -9234 -33633 -9198
rect -33417 -9243 -33390 -9216
rect -33867 -9279 -33849 -9261
rect -33417 -9261 -33318 -9243
rect -33417 -9279 -33381 -9261
rect -33975 -9297 -33381 -9279
rect -35388 -9396 -35370 -9369
rect -34335 -9423 -34317 -9414
rect -33975 -9810 -33957 -9297
rect -33678 -9360 -33660 -9351
rect -33192 -9513 -33174 -9000
rect -31437 -9126 -31419 -9117
rect -31284 -9468 -31266 -9414
rect -33417 -9531 -33174 -9513
rect -33417 -9558 -33390 -9531
rect -33867 -9576 -33390 -9558
rect -33867 -9630 -33849 -9576
rect -33714 -9630 -33696 -9576
rect -33417 -9585 -33390 -9576
rect -33813 -9711 -33795 -9657
rect -33651 -9711 -33633 -9648
rect -33345 -9666 -33318 -9621
rect -33489 -9702 -33399 -9675
rect -33345 -9693 -33327 -9666
rect -33489 -9711 -33471 -9702
rect -33813 -9729 -33471 -9711
rect -33345 -9711 -33318 -9693
rect -33651 -9765 -33633 -9729
rect -33417 -9774 -33390 -9747
rect -33867 -9810 -33849 -9792
rect -33417 -9792 -33318 -9774
rect -33417 -9810 -33381 -9792
rect -33975 -9828 -33381 -9810
rect -35298 -9954 -35289 -9936
rect -35271 -9954 -35253 -9936
rect -34452 -9990 -34434 -9963
rect -33975 -10287 -33957 -9828
rect -33678 -9927 -33660 -9891
rect -33192 -9990 -33174 -9531
rect -31392 -9693 -31374 -9666
rect -33417 -10008 -33174 -9990
rect -33417 -10035 -33390 -10008
rect -33867 -10053 -33390 -10035
rect -33867 -10107 -33849 -10053
rect -33714 -10107 -33696 -10053
rect -33417 -10062 -33390 -10053
rect -33813 -10188 -33795 -10134
rect -33651 -10188 -33633 -10125
rect -33345 -10143 -33318 -10098
rect -33489 -10179 -33399 -10152
rect -33345 -10170 -33327 -10143
rect -33489 -10188 -33471 -10179
rect -33813 -10206 -33471 -10188
rect -33345 -10188 -33318 -10170
rect -33651 -10242 -33633 -10206
rect -33417 -10251 -33390 -10224
rect -33867 -10287 -33849 -10269
rect -33417 -10269 -33318 -10251
rect -33417 -10287 -33381 -10269
rect -33975 -10305 -33381 -10287
rect -34614 -10413 -34578 -10395
rect -33975 -10782 -33957 -10305
rect -33678 -10386 -33660 -10359
rect -33192 -10485 -33174 -10008
rect -31230 -10413 -31212 -8748
rect -30960 -10341 -30942 -5634
rect -30879 -7020 -30861 -6813
rect -30960 -10377 -30942 -10368
rect -30843 -9423 -30825 -5571
rect -30402 -5553 -29520 -5535
rect -30402 -6246 -30384 -5553
rect -29340 -5760 -29322 -5004
rect -29160 -5049 -29133 -5004
rect -28827 -5058 -28809 -5004
rect -28674 -5058 -28656 -5004
rect -28377 -5013 -28350 -5004
rect -29169 -5166 -29160 -5139
rect -29088 -5175 -29061 -5085
rect -28773 -5139 -28755 -5085
rect -28611 -5139 -28593 -5076
rect -28449 -5130 -28359 -5103
rect -28449 -5139 -28431 -5130
rect -28773 -5157 -28431 -5139
rect -28305 -5139 -28278 -5049
rect -27999 -5058 -27981 -5004
rect -27846 -5058 -27828 -5004
rect -27549 -5013 -27522 -5004
rect -27126 -5013 -27108 -4959
rect -28611 -5193 -28593 -5157
rect -29160 -5238 -29133 -5211
rect -27945 -5139 -27927 -5085
rect -27783 -5139 -27765 -5076
rect -27477 -5094 -27450 -5049
rect -27126 -5031 -26676 -5013
rect -27126 -5067 -27108 -5031
rect -26721 -5067 -26703 -5031
rect -27621 -5130 -27531 -5103
rect -27477 -5121 -27270 -5094
rect -27621 -5139 -27603 -5130
rect -27945 -5157 -27603 -5139
rect -27477 -5139 -27450 -5121
rect -28377 -5202 -28350 -5175
rect -27783 -5193 -27765 -5157
rect -28827 -5238 -28809 -5220
rect -28377 -5220 -28278 -5202
rect -27288 -5130 -27270 -5121
rect -27288 -5148 -27090 -5130
rect -26793 -5148 -26775 -5094
rect -26667 -5148 -26649 -5094
rect -27063 -5166 -26694 -5148
rect -26667 -5166 -26622 -5148
rect -27549 -5202 -27522 -5175
rect -27063 -5193 -27045 -5166
rect -26973 -5193 -26955 -5166
rect -26883 -5193 -26865 -5166
rect -26793 -5193 -26775 -5166
rect -26667 -5193 -26649 -5166
rect -28377 -5238 -28341 -5220
rect -27999 -5238 -27981 -5220
rect -27549 -5220 -27450 -5202
rect -27549 -5238 -27513 -5220
rect -27126 -5238 -27108 -5211
rect -27027 -5238 -27009 -5211
rect -26937 -5238 -26919 -5211
rect -26847 -5238 -26829 -5211
rect -26721 -5238 -26703 -5211
rect -29124 -5256 -26703 -5238
rect -29340 -5787 -27846 -5760
rect -30078 -5832 -29862 -5796
rect -29826 -5832 -29646 -5796
rect -29340 -5823 -29322 -5787
rect -30078 -5904 -29862 -5868
rect -29826 -5904 -29691 -5868
rect -30240 -6003 -30114 -5967
rect -30078 -6003 -29862 -5967
rect -29727 -5985 -29691 -5904
rect -30240 -6102 -30204 -6003
rect -29727 -6021 -29718 -5985
rect -29727 -6039 -29691 -6021
rect -30078 -6075 -29862 -6039
rect -29826 -6075 -29691 -6039
rect -29682 -6102 -29646 -5832
rect -30240 -6138 -30015 -6102
rect -30240 -6192 -30114 -6156
rect -30240 -6246 -30204 -6228
rect -30051 -6237 -30015 -6138
rect -29997 -6138 -29646 -6102
rect -29610 -5832 -29322 -5823
rect -28674 -5832 -28647 -5787
rect -29610 -5841 -29079 -5832
rect -29997 -6147 -29961 -6138
rect -29826 -6192 -29709 -6156
rect -30402 -6264 -30204 -6246
rect -30402 -6552 -30384 -6264
rect -30240 -6282 -30204 -6264
rect -30078 -6273 -29862 -6237
rect -29745 -6246 -29709 -6228
rect -29610 -6246 -29583 -5841
rect -29520 -5850 -29484 -5841
rect -29511 -5895 -29484 -5850
rect -29340 -5850 -29151 -5841
rect -29439 -6021 -29412 -5931
rect -29511 -6084 -29484 -6057
rect -29745 -6273 -29583 -6246
rect -29538 -6102 -29457 -6084
rect -29745 -6282 -29709 -6273
rect -30240 -6354 -30114 -6318
rect -29943 -6327 -29925 -6309
rect -29826 -6354 -29709 -6318
rect -30240 -6408 -30222 -6390
rect -30078 -6435 -29862 -6399
rect -29997 -6462 -29961 -6435
rect -29943 -6498 -29925 -6480
rect -29538 -6552 -29520 -6102
rect -30402 -6570 -29520 -6552
rect -30402 -7542 -30384 -6570
rect -29340 -7056 -29322 -5850
rect -29178 -5895 -29151 -5850
rect -28548 -5832 -28521 -5787
rect -28404 -5832 -28377 -5787
rect -28611 -5913 -28584 -5868
rect -28278 -5832 -28251 -5787
rect -28485 -5913 -28458 -5868
rect -28152 -5832 -28125 -5787
rect -28341 -5913 -28314 -5868
rect -27882 -5823 -27855 -5787
rect -28215 -5913 -28188 -5868
rect -28080 -5913 -28053 -5868
rect -27819 -5913 -27792 -5868
rect -26946 -5913 -26928 -5562
rect -29106 -5976 -29079 -5931
rect -28881 -5958 -28656 -5931
rect -28611 -5940 -27855 -5913
rect -27819 -5940 -26928 -5913
rect -28881 -5976 -28863 -5958
rect -28278 -5976 -28251 -5949
rect -29106 -6003 -28863 -5976
rect -28053 -6003 -28026 -5940
rect -27819 -6003 -27792 -5940
rect -29106 -6021 -29079 -6003
rect -29178 -6084 -29151 -6057
rect -28674 -6075 -28647 -6030
rect -27882 -6075 -27855 -6030
rect -28674 -6084 -27855 -6075
rect -29187 -6102 -29178 -6084
rect -29142 -6102 -27855 -6084
rect -29340 -7065 -27999 -7056
rect -30078 -7128 -29862 -7092
rect -29826 -7128 -29646 -7092
rect -30078 -7200 -29862 -7164
rect -29826 -7200 -29691 -7164
rect -30240 -7299 -30114 -7263
rect -30078 -7299 -29862 -7263
rect -29727 -7281 -29691 -7200
rect -30240 -7398 -30204 -7299
rect -29727 -7317 -29718 -7281
rect -29727 -7335 -29691 -7317
rect -30078 -7371 -29862 -7335
rect -29826 -7371 -29691 -7335
rect -29682 -7398 -29646 -7128
rect -30240 -7434 -30015 -7398
rect -30240 -7488 -30114 -7452
rect -30240 -7542 -30204 -7524
rect -30051 -7533 -30015 -7434
rect -29997 -7434 -29646 -7398
rect -29610 -7137 -29340 -7119
rect -29322 -7083 -27999 -7065
rect -29322 -7137 -29133 -7119
rect -28827 -7128 -28800 -7083
rect -29997 -7443 -29961 -7434
rect -29826 -7488 -29709 -7452
rect -30402 -7560 -30204 -7542
rect -30402 -7848 -30384 -7560
rect -30240 -7578 -30204 -7560
rect -30078 -7569 -29862 -7533
rect -29745 -7542 -29709 -7524
rect -29610 -7542 -29583 -7137
rect -29520 -7146 -29484 -7137
rect -29241 -7146 -29205 -7137
rect -29511 -7191 -29484 -7146
rect -29232 -7191 -29205 -7146
rect -28701 -7128 -28674 -7083
rect -28557 -7128 -28530 -7083
rect -29439 -7272 -29412 -7227
rect -28764 -7209 -28737 -7164
rect -28431 -7128 -28404 -7083
rect -28638 -7209 -28611 -7164
rect -28305 -7128 -28278 -7083
rect -28494 -7209 -28467 -7164
rect -28035 -7119 -28008 -7083
rect -28368 -7209 -28341 -7164
rect -28233 -7209 -28206 -7164
rect -27972 -7209 -27945 -7164
rect -26856 -7209 -26838 -5976
rect -29160 -7272 -29133 -7227
rect -28971 -7254 -28809 -7227
rect -28764 -7236 -28008 -7209
rect -27972 -7236 -26838 -7209
rect -28971 -7272 -28953 -7254
rect -29439 -7299 -29385 -7272
rect -29439 -7317 -29412 -7299
rect -29160 -7299 -28953 -7272
rect -28206 -7299 -28179 -7236
rect -27972 -7299 -27945 -7236
rect -29160 -7317 -29133 -7299
rect -29511 -7380 -29484 -7353
rect -29232 -7380 -29205 -7353
rect -28827 -7371 -28800 -7326
rect -28035 -7371 -28008 -7326
rect -28827 -7380 -28008 -7371
rect -29745 -7569 -29583 -7542
rect -29538 -7398 -28008 -7380
rect -29745 -7578 -29709 -7569
rect -29943 -7614 -29925 -7605
rect -30240 -7650 -30114 -7614
rect -29826 -7650 -29709 -7614
rect -30078 -7731 -29862 -7695
rect -29997 -7758 -29961 -7731
rect -29538 -7848 -29520 -7398
rect -30402 -7866 -29520 -7848
rect -30402 -9081 -30384 -7866
rect -30078 -8667 -29862 -8631
rect -29826 -8667 -29646 -8631
rect -30078 -8739 -29862 -8703
rect -29826 -8739 -29691 -8703
rect -30240 -8838 -30114 -8802
rect -30078 -8838 -29862 -8802
rect -29727 -8820 -29691 -8739
rect -30240 -8937 -30204 -8838
rect -29727 -8856 -29718 -8820
rect -29727 -8874 -29691 -8856
rect -30078 -8910 -29862 -8874
rect -29826 -8910 -29691 -8874
rect -29682 -8937 -29646 -8667
rect -30240 -8973 -30015 -8937
rect -30240 -9027 -30114 -8991
rect -30240 -9081 -30204 -9063
rect -30402 -9099 -30204 -9081
rect -30402 -9387 -30384 -9099
rect -30240 -9117 -30204 -9099
rect -30186 -9081 -30168 -9063
rect -30051 -9072 -30015 -8973
rect -29997 -8973 -29646 -8937
rect -29610 -8676 -29340 -8658
rect -29997 -8982 -29961 -8973
rect -29826 -9027 -29709 -8991
rect -30078 -9108 -29862 -9072
rect -29745 -9081 -29709 -9063
rect -29610 -9081 -29583 -8676
rect -29520 -8685 -29484 -8676
rect -29511 -8730 -29484 -8685
rect -29439 -8856 -29412 -8766
rect -29511 -8919 -29484 -8892
rect -29745 -9108 -29583 -9081
rect -29538 -8937 -29421 -8919
rect -29745 -9117 -29709 -9108
rect -30240 -9189 -30114 -9153
rect -29826 -9189 -29709 -9153
rect -30078 -9270 -29862 -9234
rect -29997 -9297 -29961 -9270
rect -29538 -9387 -29520 -8937
rect -30402 -9405 -29520 -9387
rect -30843 -10449 -30825 -9441
rect -31383 -10467 -30825 -10449
rect -30402 -10026 -30384 -9405
rect -29781 -9468 -29763 -9450
rect -30078 -9612 -29862 -9576
rect -29826 -9612 -29646 -9576
rect -29340 -9603 -29322 -8721
rect -30078 -9684 -29862 -9648
rect -29826 -9684 -29691 -9648
rect -30240 -9783 -30114 -9747
rect -30078 -9783 -29862 -9747
rect -29727 -9765 -29691 -9684
rect -30240 -9882 -30204 -9783
rect -29727 -9801 -29718 -9765
rect -29727 -9819 -29691 -9801
rect -30078 -9855 -29862 -9819
rect -29826 -9855 -29691 -9819
rect -29682 -9882 -29646 -9612
rect -30240 -9918 -30015 -9882
rect -30240 -9972 -30114 -9936
rect -30240 -10026 -30204 -10008
rect -30402 -10044 -30204 -10026
rect -30402 -10332 -30384 -10044
rect -30240 -10062 -30204 -10044
rect -30186 -10026 -30168 -10008
rect -30051 -10017 -30015 -9918
rect -29997 -9918 -29646 -9882
rect -29610 -9621 -28179 -9603
rect -29997 -9927 -29961 -9918
rect -29826 -9972 -29709 -9936
rect -30078 -10053 -29862 -10017
rect -29745 -10026 -29709 -10008
rect -29610 -10026 -29583 -9621
rect -29520 -9630 -29484 -9621
rect -29511 -9675 -29484 -9630
rect -29439 -9801 -29412 -9711
rect -29511 -9864 -29484 -9837
rect -29745 -10053 -29583 -10026
rect -29538 -9882 -29421 -9864
rect -29745 -10062 -29709 -10053
rect -30240 -10134 -30114 -10098
rect -29826 -10134 -29709 -10098
rect -30078 -10215 -29862 -10179
rect -29997 -10242 -29961 -10215
rect -29538 -10332 -29520 -9882
rect -30402 -10350 -29556 -10332
rect -33417 -10503 -33174 -10485
rect -33417 -10530 -33390 -10503
rect -33867 -10548 -33390 -10530
rect -33867 -10602 -33849 -10548
rect -33714 -10602 -33696 -10548
rect -33417 -10557 -33390 -10548
rect -33813 -10683 -33795 -10629
rect -33651 -10683 -33633 -10620
rect -33345 -10638 -33318 -10593
rect -33489 -10674 -33399 -10647
rect -33345 -10665 -33327 -10638
rect -33489 -10683 -33471 -10674
rect -33813 -10701 -33471 -10683
rect -33345 -10683 -33318 -10665
rect -33651 -10737 -33633 -10701
rect -33417 -10746 -33390 -10719
rect -33867 -10782 -33849 -10764
rect -33417 -10764 -33318 -10746
rect -33417 -10782 -33381 -10764
rect -33975 -10800 -33381 -10782
rect -34776 -10881 -34740 -10863
rect -33975 -11196 -33957 -10800
rect -33678 -10863 -33660 -10854
rect -33192 -10899 -33174 -10503
rect -31473 -10665 -30960 -10638
rect -33417 -10917 -33174 -10899
rect -33417 -10944 -33390 -10917
rect -33867 -10962 -33390 -10944
rect -33867 -11016 -33849 -10962
rect -33714 -11016 -33696 -10962
rect -33417 -10971 -33390 -10962
rect -33813 -11097 -33795 -11043
rect -33651 -11097 -33633 -11034
rect -33345 -11052 -33318 -11007
rect -33489 -11088 -33399 -11061
rect -33345 -11079 -33327 -11052
rect -33489 -11097 -33471 -11088
rect -33813 -11115 -33471 -11097
rect -33345 -11097 -33318 -11079
rect -33651 -11151 -33633 -11115
rect -33417 -11160 -33390 -11133
rect -33867 -11196 -33849 -11178
rect -33417 -11178 -33318 -11160
rect -33417 -11196 -33381 -11178
rect -33975 -11214 -33381 -11196
rect -36207 -11313 -35217 -11295
rect -36207 -12078 -36189 -11313
rect -35244 -11412 -35217 -11313
rect -34947 -11313 -34920 -11295
rect -35415 -11430 -35217 -11412
rect -35415 -11457 -35388 -11430
rect -35865 -11475 -35388 -11457
rect -35865 -11529 -35847 -11475
rect -35712 -11529 -35694 -11475
rect -35415 -11484 -35388 -11475
rect -35811 -11610 -35793 -11556
rect -35649 -11610 -35631 -11547
rect -35343 -11565 -35316 -11520
rect -35487 -11601 -35397 -11574
rect -35343 -11592 -35325 -11565
rect -35487 -11610 -35469 -11601
rect -35865 -11637 -35847 -11619
rect -35811 -11628 -35469 -11610
rect -35343 -11610 -35316 -11592
rect -35712 -11655 -35694 -11637
rect -35649 -11664 -35631 -11628
rect -35415 -11673 -35388 -11646
rect -35865 -11709 -35847 -11691
rect -35415 -11691 -35316 -11673
rect -35415 -11709 -35379 -11691
rect -35955 -11727 -35379 -11709
rect -36216 -12096 -36108 -12078
rect -36207 -12141 -36180 -12096
rect -36135 -12222 -36108 -12177
rect -35955 -12177 -35937 -11727
rect -35244 -11880 -35217 -11430
rect -33975 -11709 -33957 -11214
rect -33678 -11295 -33660 -11259
rect -33192 -11430 -33174 -10917
rect -33417 -11448 -33174 -11430
rect -33417 -11475 -33390 -11448
rect -33867 -11493 -33390 -11475
rect -33867 -11547 -33849 -11493
rect -33714 -11547 -33696 -11493
rect -33417 -11502 -33390 -11493
rect -33813 -11628 -33795 -11574
rect -33651 -11628 -33633 -11565
rect -33345 -11583 -33318 -11538
rect -33489 -11619 -33399 -11592
rect -33345 -11610 -33336 -11583
rect -33489 -11628 -33471 -11619
rect -33813 -11646 -33471 -11628
rect -33345 -11628 -33318 -11610
rect -33651 -11682 -33633 -11646
rect -33417 -11691 -33390 -11664
rect -33192 -11682 -33174 -11448
rect -30402 -11043 -30384 -10350
rect -29781 -10413 -29763 -10404
rect -30078 -10629 -29862 -10593
rect -29826 -10629 -29646 -10593
rect -29340 -10620 -29322 -9621
rect -28206 -9711 -28179 -9621
rect -26406 -9684 -26307 -9675
rect -26406 -9711 -26379 -9684
rect -28206 -9729 -26379 -9711
rect -28206 -9738 -27378 -9729
rect -28206 -9783 -28179 -9738
rect -28080 -9783 -28053 -9738
rect -27936 -9783 -27909 -9738
rect -28143 -9864 -28116 -9819
rect -27810 -9783 -27783 -9738
rect -28017 -9864 -27990 -9819
rect -27684 -9783 -27657 -9738
rect -27873 -9864 -27846 -9819
rect -27414 -9774 -27387 -9738
rect -27747 -9864 -27720 -9819
rect -26856 -9783 -26838 -9729
rect -27612 -9864 -27585 -9819
rect -26703 -9783 -26685 -9729
rect -26406 -9738 -26379 -9729
rect -28143 -9891 -27387 -9864
rect -27585 -9954 -27558 -9891
rect -27351 -9954 -27324 -9819
rect -26802 -9864 -26784 -9810
rect -26640 -9864 -26622 -9801
rect -26334 -9819 -26307 -9774
rect -26478 -9855 -26388 -9828
rect -26334 -9846 -26280 -9819
rect -26478 -9864 -26460 -9855
rect -26802 -9882 -26460 -9864
rect -26334 -9864 -26307 -9846
rect -26640 -9918 -26622 -9882
rect -26406 -9927 -26379 -9900
rect -26856 -9963 -26838 -9945
rect -26406 -9945 -26307 -9927
rect -26406 -9963 -26370 -9945
rect -26856 -9981 -26370 -9963
rect -28206 -10026 -28179 -9981
rect -27414 -10026 -27387 -9981
rect -26838 -10026 -26820 -9981
rect -28206 -10053 -26820 -10026
rect -28188 -10314 -28170 -10053
rect -30078 -10701 -29862 -10665
rect -29826 -10701 -29691 -10665
rect -30240 -10800 -30114 -10764
rect -30078 -10800 -29862 -10764
rect -29727 -10782 -29691 -10701
rect -30240 -10899 -30204 -10800
rect -29727 -10818 -29718 -10782
rect -29727 -10836 -29691 -10818
rect -30078 -10872 -29862 -10836
rect -29826 -10872 -29691 -10836
rect -29682 -10899 -29646 -10629
rect -30240 -10935 -30015 -10899
rect -30240 -10989 -30114 -10953
rect -30240 -11043 -30204 -11025
rect -30051 -11034 -30015 -10935
rect -29997 -10935 -29646 -10899
rect -29610 -10638 -29322 -10620
rect -29997 -10944 -29961 -10935
rect -29826 -10989 -29709 -10953
rect -30402 -11061 -30204 -11043
rect -30402 -11349 -30384 -11061
rect -30240 -11079 -30204 -11061
rect -30078 -11070 -29862 -11034
rect -29745 -11043 -29709 -11025
rect -29610 -11043 -29583 -10638
rect -29520 -10647 -29484 -10638
rect -29511 -10692 -29484 -10647
rect -29439 -10818 -29412 -10728
rect -29511 -10881 -29484 -10854
rect -29745 -11070 -29583 -11043
rect -29538 -10899 -29421 -10881
rect -29745 -11079 -29709 -11070
rect -30240 -11151 -30114 -11115
rect -29826 -11151 -29709 -11115
rect -30339 -11187 -30285 -11169
rect -30078 -11232 -29862 -11196
rect -29997 -11259 -29961 -11232
rect -29538 -11349 -29520 -10899
rect -30402 -11367 -29520 -11349
rect -31203 -11610 -31176 -11583
rect -33867 -11727 -33849 -11709
rect -33417 -11709 -33318 -11691
rect -33417 -11727 -33381 -11709
rect -33957 -11745 -33381 -11727
rect -33678 -11871 -33660 -11826
rect -35415 -11898 -35217 -11880
rect -35415 -11925 -35388 -11898
rect -35865 -11943 -35388 -11925
rect -35865 -11997 -35847 -11943
rect -35712 -11997 -35694 -11943
rect -35415 -11952 -35388 -11943
rect -35811 -12078 -35793 -12024
rect -35649 -12078 -35631 -12015
rect -35343 -12033 -35316 -11988
rect -35487 -12069 -35397 -12042
rect -35343 -12060 -35334 -12033
rect -35487 -12078 -35469 -12069
rect -35811 -12096 -35469 -12078
rect -35343 -12078 -35316 -12060
rect -35703 -12123 -35676 -12105
rect -35649 -12132 -35631 -12096
rect -35415 -12141 -35388 -12114
rect -35865 -12177 -35847 -12159
rect -35415 -12159 -35316 -12141
rect -35415 -12177 -35379 -12159
rect -35955 -12195 -35379 -12177
rect -36135 -12249 -36054 -12222
rect -36135 -12267 -36108 -12249
rect -36207 -12330 -36180 -12303
rect -35955 -12330 -35937 -12195
rect -35244 -12321 -35217 -11898
rect -35127 -11898 -35100 -11880
rect -33192 -12294 -33174 -11718
rect -36333 -12348 -35937 -12330
rect -35415 -12339 -35217 -12321
rect -33417 -12312 -33174 -12294
rect -33417 -12339 -33390 -12312
rect -36333 -12654 -36315 -12348
rect -35415 -12366 -35388 -12339
rect -35973 -12384 -35388 -12366
rect -35973 -12393 -35955 -12384
rect -36207 -12411 -35955 -12393
rect -36207 -12420 -36171 -12411
rect -36198 -12465 -36171 -12420
rect -35865 -12438 -35847 -12384
rect -35712 -12438 -35694 -12384
rect -35415 -12393 -35388 -12384
rect -35244 -12357 -33390 -12339
rect -36126 -12546 -36099 -12501
rect -35811 -12519 -35793 -12465
rect -35649 -12519 -35631 -12456
rect -35343 -12474 -35316 -12429
rect -35487 -12510 -35397 -12483
rect -35343 -12501 -35334 -12474
rect -35487 -12519 -35469 -12510
rect -35874 -12537 -35838 -12519
rect -35811 -12537 -35469 -12519
rect -35343 -12519 -35316 -12501
rect -36126 -12573 -36063 -12546
rect -35649 -12573 -35631 -12537
rect -36126 -12591 -36099 -12573
rect -35415 -12582 -35388 -12555
rect -35865 -12618 -35847 -12600
rect -35415 -12600 -35316 -12582
rect -35415 -12618 -35379 -12600
rect -36198 -12654 -36171 -12627
rect -35865 -12636 -35379 -12618
rect -35865 -12654 -35847 -12636
rect -36333 -12672 -35847 -12654
rect -36198 -13014 -36180 -12672
rect -35244 -12735 -35217 -12357
rect -33867 -12411 -33849 -12357
rect -33714 -12411 -33696 -12357
rect -33417 -12366 -33390 -12357
rect -33201 -12321 -33174 -12312
rect -33813 -12492 -33795 -12438
rect -33651 -12492 -33633 -12429
rect -33345 -12447 -33318 -12402
rect -33489 -12483 -33399 -12456
rect -33345 -12474 -33336 -12447
rect -33489 -12492 -33471 -12483
rect -33813 -12510 -33471 -12492
rect -33345 -12492 -33318 -12474
rect -33651 -12546 -33633 -12510
rect -33417 -12555 -33390 -12528
rect -33867 -12591 -33849 -12573
rect -33417 -12591 -33381 -12555
rect -35415 -12753 -35217 -12735
rect -33957 -12609 -33381 -12591
rect -35415 -12780 -35388 -12753
rect -35865 -12798 -35388 -12780
rect -35865 -12852 -35847 -12798
rect -35712 -12852 -35694 -12798
rect -35415 -12807 -35388 -12798
rect -35811 -12933 -35793 -12879
rect -35649 -12933 -35631 -12870
rect -35343 -12888 -35316 -12843
rect -35487 -12924 -35397 -12897
rect -35343 -12915 -35334 -12888
rect -35487 -12933 -35469 -12924
rect -35811 -12951 -35469 -12933
rect -35343 -12933 -35316 -12915
rect -35649 -12987 -35631 -12951
rect -36207 -13032 -36180 -13014
rect -35415 -12996 -35388 -12969
rect -35865 -13032 -35847 -13014
rect -35415 -13014 -35307 -12996
rect -35415 -13032 -35379 -13014
rect -36207 -13050 -35379 -13032
rect -36207 -13428 -36189 -13050
rect -35352 -13068 -35307 -13014
rect -33975 -13068 -33957 -12645
rect -33201 -12789 -33183 -12321
rect -30402 -12339 -30384 -11367
rect -29340 -11673 -29322 -10638
rect -30078 -11925 -29862 -11889
rect -29826 -11925 -29646 -11889
rect -29340 -11916 -29322 -11718
rect -30078 -11997 -29862 -11961
rect -29826 -11997 -29691 -11961
rect -30240 -12096 -30114 -12060
rect -30078 -12096 -29862 -12060
rect -29727 -12078 -29691 -11997
rect -30240 -12195 -30204 -12096
rect -29727 -12114 -29718 -12078
rect -29727 -12132 -29691 -12114
rect -30078 -12168 -29862 -12132
rect -29826 -12168 -29691 -12132
rect -29682 -12195 -29646 -11925
rect -30240 -12231 -30015 -12195
rect -30240 -12285 -30114 -12249
rect -30240 -12339 -30204 -12321
rect -30051 -12330 -30015 -12231
rect -29997 -12231 -29646 -12195
rect -29610 -11934 -29322 -11916
rect -29997 -12240 -29961 -12231
rect -29826 -12285 -29709 -12249
rect -30402 -12357 -30204 -12339
rect -30402 -12546 -30384 -12357
rect -30240 -12375 -30204 -12357
rect -30078 -12366 -29862 -12330
rect -29745 -12339 -29709 -12321
rect -29610 -12339 -29583 -11934
rect -29520 -11943 -29484 -11934
rect -29511 -11988 -29484 -11943
rect -29439 -12114 -29412 -12024
rect -29511 -12177 -29484 -12150
rect -29745 -12366 -29583 -12339
rect -29538 -12195 -29421 -12177
rect -29745 -12375 -29709 -12366
rect -30240 -12447 -30114 -12411
rect -29826 -12447 -29709 -12411
rect -30078 -12528 -29862 -12492
rect -29997 -12555 -29961 -12528
rect -30402 -12645 -30384 -12600
rect -29538 -12645 -29520 -12195
rect -30402 -12663 -29520 -12645
rect -31374 -12681 -31356 -12663
rect -33417 -12807 -33183 -12789
rect -33417 -12834 -33390 -12807
rect -33867 -12852 -33390 -12834
rect -33867 -12906 -33849 -12852
rect -33714 -12906 -33696 -12852
rect -33417 -12861 -33390 -12852
rect -33813 -12987 -33795 -12933
rect -33651 -12987 -33633 -12924
rect -33345 -12942 -33318 -12897
rect -33489 -12978 -33399 -12951
rect -33345 -12969 -33336 -12942
rect -33489 -12987 -33471 -12978
rect -33813 -13005 -33471 -12987
rect -33345 -12987 -33318 -12969
rect -33651 -13041 -33633 -13005
rect -35352 -13086 -33957 -13068
rect -33417 -13050 -33390 -13023
rect -33867 -13086 -33849 -13068
rect -33417 -13068 -33318 -13050
rect -33417 -13086 -33381 -13068
rect -37332 -13455 -36189 -13428
rect -37332 -13500 -37296 -13455
rect -36207 -13464 -36189 -13455
rect -33975 -13104 -33381 -13086
rect -33975 -13500 -33957 -13104
rect -33678 -13140 -33660 -13131
rect -33201 -13203 -33183 -12807
rect -33417 -13221 -33183 -13203
rect -33417 -13248 -33390 -13221
rect -33867 -13266 -33390 -13248
rect -33867 -13320 -33849 -13266
rect -33714 -13320 -33696 -13266
rect -33417 -13275 -33390 -13266
rect -33813 -13401 -33795 -13347
rect -33651 -13401 -33633 -13338
rect -33345 -13356 -33318 -13311
rect -33489 -13392 -33399 -13365
rect -33345 -13383 -33327 -13356
rect -33489 -13401 -33471 -13392
rect -33813 -13419 -33471 -13401
rect -33345 -13401 -33318 -13383
rect -33651 -13455 -33633 -13419
rect -33417 -13464 -33390 -13437
rect -33867 -13500 -33849 -13482
rect -33417 -13482 -33318 -13464
rect -33417 -13500 -33381 -13482
rect -33975 -13518 -33381 -13500
rect -33975 -14031 -33957 -13518
rect -33678 -13617 -33660 -13590
rect -33201 -13734 -33183 -13221
rect -33417 -13752 -33183 -13734
rect -33417 -13779 -33390 -13752
rect -33867 -13797 -33390 -13779
rect -33867 -13851 -33849 -13797
rect -33714 -13851 -33696 -13797
rect -33417 -13806 -33390 -13797
rect -33813 -13932 -33795 -13878
rect -33651 -13932 -33633 -13869
rect -33345 -13887 -33318 -13842
rect -33489 -13923 -33399 -13896
rect -33345 -13914 -33336 -13887
rect -33489 -13932 -33471 -13923
rect -33813 -13950 -33471 -13932
rect -33345 -13932 -33318 -13914
rect -33651 -13986 -33633 -13950
rect -33417 -13995 -33390 -13968
rect -33867 -14031 -33849 -14013
rect -33417 -14013 -33318 -13995
rect -33417 -14031 -33381 -14013
rect -33975 -14049 -33381 -14031
rect -33975 -14526 -33957 -14049
rect -33678 -14112 -33660 -14094
rect -33201 -14229 -33183 -13752
rect -31446 -13761 -31347 -13752
rect -31446 -13788 -31419 -13761
rect -33417 -14247 -33183 -14229
rect -33417 -14274 -33390 -14247
rect -33867 -14292 -33390 -14274
rect -33867 -14346 -33849 -14292
rect -33714 -14346 -33696 -14292
rect -33417 -14301 -33390 -14292
rect -33813 -14427 -33795 -14373
rect -33651 -14427 -33633 -14364
rect -33345 -14382 -33318 -14337
rect -33489 -14418 -33399 -14391
rect -33345 -14409 -33327 -14382
rect -33489 -14427 -33471 -14418
rect -33813 -14445 -33471 -14427
rect -33345 -14427 -33318 -14409
rect -33651 -14481 -33633 -14445
rect -33417 -14490 -33390 -14463
rect -33867 -14526 -33849 -14508
rect -33417 -14508 -33354 -14490
rect -33417 -14526 -33381 -14508
rect -33975 -14544 -33381 -14526
rect -33975 -15021 -33957 -14544
rect -33678 -14607 -33660 -14598
rect -33201 -14652 -33183 -14247
rect -32058 -13806 -31419 -13788
rect -32058 -14265 -32040 -13806
rect -31896 -13860 -31878 -13806
rect -31743 -13860 -31725 -13806
rect -31446 -13815 -31419 -13806
rect -31842 -13941 -31824 -13887
rect -31680 -13941 -31662 -13878
rect -31374 -13896 -31347 -13851
rect -31518 -13932 -31428 -13905
rect -31374 -13923 -31320 -13896
rect -31518 -13941 -31500 -13932
rect -31842 -13959 -31500 -13941
rect -31374 -13941 -31347 -13923
rect -31680 -13995 -31662 -13959
rect -31446 -14004 -31419 -13977
rect -31896 -14040 -31878 -14022
rect -31446 -14022 -31230 -14004
rect -31446 -14040 -31410 -14022
rect -31896 -14058 -31410 -14040
rect -31869 -14139 -31851 -14112
rect -31707 -14112 -31689 -14103
rect -31446 -14238 -31347 -14229
rect -31446 -14265 -31419 -14238
rect -32058 -14283 -31419 -14265
rect -32058 -14652 -32040 -14283
rect -31896 -14337 -31878 -14283
rect -31743 -14337 -31725 -14283
rect -31446 -14292 -31419 -14283
rect -31842 -14418 -31824 -14364
rect -31680 -14418 -31662 -14355
rect -31374 -14373 -31347 -14328
rect -31518 -14409 -31428 -14382
rect -31374 -14400 -31320 -14373
rect -31518 -14418 -31500 -14409
rect -31842 -14436 -31500 -14418
rect -31374 -14418 -31347 -14400
rect -31680 -14472 -31662 -14436
rect -31446 -14481 -31419 -14454
rect -31248 -14481 -31230 -14022
rect -31896 -14517 -31878 -14499
rect -31446 -14499 -31230 -14481
rect -31446 -14517 -31410 -14499
rect -31896 -14535 -31410 -14517
rect -31869 -14616 -31851 -14571
rect -31707 -14589 -31689 -14580
rect -31446 -14634 -31347 -14625
rect -33201 -14661 -32040 -14652
rect -31446 -14661 -31419 -14634
rect -33201 -14679 -31419 -14661
rect -33201 -14688 -32040 -14679
rect -33201 -14724 -33183 -14688
rect -33417 -14742 -33183 -14724
rect -33417 -14769 -33390 -14742
rect -33867 -14787 -33390 -14769
rect -33867 -14841 -33849 -14787
rect -33714 -14841 -33696 -14787
rect -33417 -14796 -33390 -14787
rect -33813 -14922 -33795 -14868
rect -33651 -14922 -33633 -14859
rect -33345 -14877 -33318 -14832
rect -33489 -14913 -33399 -14886
rect -33345 -14904 -33327 -14877
rect -33489 -14922 -33471 -14913
rect -33813 -14940 -33471 -14922
rect -33345 -14922 -33318 -14904
rect -33651 -14976 -33633 -14940
rect -33417 -14985 -33390 -14958
rect -33867 -15021 -33849 -15003
rect -33417 -15003 -33318 -14985
rect -33417 -15021 -33381 -15003
rect -33975 -15039 -33381 -15021
rect -33975 -15435 -33957 -15039
rect -33678 -15093 -33660 -15075
rect -33201 -15138 -33183 -14742
rect -33417 -15156 -33183 -15138
rect -32058 -15129 -32040 -14688
rect -31896 -14733 -31878 -14679
rect -31743 -14733 -31725 -14679
rect -31446 -14688 -31419 -14679
rect -31842 -14814 -31824 -14760
rect -31680 -14814 -31662 -14751
rect -31374 -14769 -31347 -14724
rect -31518 -14805 -31428 -14778
rect -31374 -14796 -31320 -14769
rect -31518 -14814 -31500 -14805
rect -31842 -14832 -31500 -14814
rect -31374 -14814 -31347 -14796
rect -31680 -14868 -31662 -14832
rect -31446 -14877 -31419 -14850
rect -31248 -14877 -31230 -14499
rect -31896 -14913 -31878 -14895
rect -31446 -14895 -31230 -14877
rect -31446 -14913 -31410 -14895
rect -31896 -14931 -31410 -14913
rect -31869 -14976 -31851 -14967
rect -31707 -15012 -31689 -15003
rect -31446 -15102 -31347 -15093
rect -31446 -15129 -31419 -15102
rect -32058 -15147 -31419 -15129
rect -33417 -15183 -33390 -15156
rect -33867 -15201 -33390 -15183
rect -33867 -15255 -33849 -15201
rect -33714 -15255 -33696 -15201
rect -33417 -15210 -33390 -15201
rect -33813 -15336 -33795 -15282
rect -33651 -15336 -33633 -15273
rect -33345 -15291 -33318 -15246
rect -33489 -15327 -33399 -15300
rect -33345 -15318 -33336 -15291
rect -33489 -15336 -33471 -15327
rect -33813 -15354 -33471 -15336
rect -33345 -15336 -33318 -15318
rect -33651 -15390 -33633 -15354
rect -33417 -15399 -33390 -15372
rect -33867 -15435 -33849 -15417
rect -33417 -15417 -33318 -15399
rect -33417 -15435 -33381 -15417
rect -33975 -15453 -33381 -15435
rect -33975 -15966 -33957 -15453
rect -33678 -15525 -33660 -15516
rect -33201 -15669 -33183 -15156
rect -31896 -15201 -31878 -15147
rect -31743 -15201 -31725 -15147
rect -31446 -15156 -31419 -15147
rect -31842 -15282 -31824 -15228
rect -31680 -15282 -31662 -15219
rect -31374 -15237 -31347 -15192
rect -31518 -15273 -31428 -15246
rect -31374 -15264 -31320 -15237
rect -31518 -15282 -31500 -15273
rect -31842 -15300 -31500 -15282
rect -31374 -15282 -31347 -15264
rect -31680 -15336 -31662 -15300
rect -33417 -15687 -33183 -15669
rect -31446 -15345 -31419 -15318
rect -31248 -15345 -31230 -14895
rect -31896 -15381 -31878 -15363
rect -31446 -15363 -31230 -15345
rect -31446 -15381 -31410 -15363
rect -31896 -15399 -31410 -15381
rect -33417 -15714 -33390 -15687
rect -33867 -15732 -33390 -15714
rect -33867 -15786 -33849 -15732
rect -33714 -15786 -33696 -15732
rect -33417 -15741 -33390 -15732
rect -33813 -15867 -33795 -15813
rect -33651 -15867 -33633 -15804
rect -33345 -15822 -33318 -15777
rect -33489 -15858 -33399 -15831
rect -33345 -15849 -33336 -15822
rect -33489 -15867 -33471 -15858
rect -33813 -15885 -33471 -15867
rect -33345 -15867 -33318 -15849
rect -33651 -15921 -33633 -15885
rect -33417 -15930 -33390 -15903
rect -31896 -15930 -31878 -15399
rect -31869 -15480 -31851 -15471
rect -31707 -15489 -31689 -15480
rect -33867 -15966 -33849 -15948
rect -33417 -15948 -31878 -15930
rect -33417 -15966 -33381 -15948
rect -33975 -15984 -33381 -15966
rect -33678 -16056 -33660 -16047
<< m2contact >>
rect -29619 10467 -29574 10485
rect -30798 9882 -30762 9900
rect -30537 9873 -30519 9900
rect -29898 9864 -29871 9891
rect -29718 9855 -29691 9891
rect -29043 9846 -29007 9882
rect -28836 9855 -28800 9882
rect -28386 9864 -28332 9882
rect -28656 9738 -28638 9765
rect -28566 9639 -28530 9657
rect -29583 8370 -29547 8388
rect -30816 7785 -30780 7803
rect -30555 7785 -30528 7803
rect -29898 7767 -29871 7794
rect -29718 7758 -29691 7794
rect -29043 7749 -29007 7785
rect -28836 7758 -28800 7785
rect -28386 7767 -28341 7785
rect -28656 7641 -28638 7668
rect -28566 7551 -28539 7569
rect -29637 6228 -29565 6264
rect -30816 5670 -30789 5688
rect -30555 5670 -30528 5688
rect -29898 5652 -29871 5679
rect -29718 5643 -29691 5679
rect -29043 5634 -29007 5670
rect -28836 5643 -28800 5670
rect -28368 5652 -28332 5670
rect -28656 5535 -28638 5562
rect -28008 5436 -27972 5454
rect -29610 4365 -29574 4383
rect -30834 3807 -30780 3825
rect -30726 3735 -30699 3744
rect -30555 3735 -30537 3744
rect -29898 3717 -29871 3744
rect -29718 3708 -29691 3744
rect -29043 3699 -29007 3735
rect -28836 3708 -28800 3735
rect -28368 3717 -28332 3735
rect -28656 3609 -28638 3627
rect -30195 63 -30168 81
rect -30843 -108 -30825 -81
rect -33354 -396 -33309 -369
rect -29943 -27 -29925 -9
rect -33354 -891 -33309 -864
rect -33354 -1305 -33309 -1278
rect -35352 -1557 -35307 -1539
rect -33705 -1566 -33669 -1530
rect -33354 -1836 -33309 -1809
rect -35235 -2115 -35181 -2079
rect -33705 -2115 -33669 -2079
rect -34596 -2655 -34551 -2628
rect -33696 -2655 -33678 -2628
rect -34758 -3123 -34713 -3087
rect -33696 -3123 -33678 -3087
rect -34947 -3627 -34893 -3600
rect -33696 -3591 -33678 -3537
rect -30717 -882 -30672 -864
rect -33345 -3843 -33309 -3816
rect -35064 -4140 -35001 -4104
rect -33696 -4095 -33678 -4050
rect -31806 -3843 -31716 -3816
rect -29151 -27 -29124 0
rect -30195 -882 -30168 -864
rect -29943 -972 -29916 -954
rect -29160 -837 -29142 -810
rect -26946 -810 -26919 -792
rect -26838 -810 -26820 -792
rect -26946 -1233 -26928 -1188
rect -31284 -6606 -31266 -6579
rect -31311 -6813 -31266 -6786
rect -35685 -8487 -35649 -8451
rect -34254 -8478 -34173 -8460
rect -35532 -8964 -35496 -8928
rect -34245 -8964 -34209 -8919
rect -33687 -8964 -33651 -8928
rect -29943 -2034 -29925 -1998
rect -29988 -2052 -29970 -2034
rect -29916 -2151 -29898 -2133
rect -28548 -1647 -28521 -1620
rect -29178 -1683 -29160 -1656
rect -26856 -1647 -26838 -1593
rect -29241 -2979 -29214 -2952
rect -29943 -3330 -29925 -3285
rect -30762 -3663 -30735 -3645
rect -30798 -3744 -30753 -3726
rect -29790 -3672 -29772 -3636
rect -29943 -4356 -29925 -4338
rect -30915 -4680 -30879 -4662
rect -29151 -4356 -29124 -4329
rect -29943 -5301 -29916 -5283
rect -30960 -5634 -30942 -5616
rect -31167 -8010 -31149 -7965
rect -35397 -9414 -35370 -9396
rect -34335 -9414 -34308 -9387
rect -33678 -9396 -33660 -9360
rect -35253 -9963 -35199 -9927
rect -34461 -9963 -34416 -9918
rect -33687 -9963 -33642 -9927
rect -34578 -10413 -34542 -10395
rect -33687 -10422 -33651 -10386
rect -30843 -5571 -30825 -5544
rect -30879 -6813 -30861 -6786
rect -30960 -10395 -30942 -10377
rect -29160 -5166 -29142 -5139
rect -26946 -5139 -26919 -5121
rect -26838 -5139 -26820 -5121
rect -26946 -5562 -26928 -5517
rect -29943 -6363 -29925 -6327
rect -29988 -6381 -29970 -6363
rect -30240 -6444 -30222 -6408
rect -29943 -6480 -29925 -6444
rect -28548 -5976 -28521 -5949
rect -29178 -6012 -29160 -5985
rect -26856 -5976 -26838 -5922
rect -29241 -7308 -29214 -7281
rect -29943 -7659 -29925 -7614
rect -30186 -9108 -30168 -9081
rect -30843 -9441 -30780 -9423
rect -30186 -10053 -30168 -10026
rect -34740 -10890 -34686 -10863
rect -33687 -10890 -33651 -10863
rect -34920 -11313 -34875 -11295
rect -35910 -11637 -35865 -11619
rect -33687 -11322 -33651 -11295
rect -31176 -11628 -31149 -11574
rect -36054 -12249 -36027 -12222
rect -35100 -11898 -35019 -11880
rect -33678 -11907 -33651 -11871
rect -35910 -12537 -35874 -12519
rect -30195 -12321 -30168 -12303
rect -33327 -14409 -33291 -14382
rect -31707 -14139 -31689 -14112
rect -31707 -14607 -31689 -14589
rect -33327 -14904 -33291 -14877
rect -31707 -15039 -31689 -15012
rect -33336 -15318 -33291 -15291
rect -33336 -15849 -33291 -15822
rect -31707 -15534 -31689 -15489
<< metal2 >>
rect -32490 10485 -32472 10494
rect -32490 10467 -29619 10485
rect -32490 -369 -32472 10467
rect -30762 9882 -30537 9900
rect -29871 9864 -29718 9882
rect -29007 9855 -28836 9882
rect -28332 9864 -27864 9882
rect -28656 9765 -28638 9774
rect -28656 9720 -28638 9738
rect -28656 9702 -28566 9720
rect -28584 9639 -28566 9702
rect -33309 -396 -32472 -369
rect -32364 8370 -29583 8388
rect -32364 -864 -32346 8370
rect -30780 7785 -30555 7803
rect -29871 7767 -29718 7785
rect -27882 7785 -27864 9864
rect -29007 7758 -28836 7785
rect -28341 7767 -27864 7785
rect -28656 7623 -28638 7641
rect -28656 7605 -28566 7623
rect -28584 7551 -28566 7605
rect -33309 -891 -32346 -864
rect -32220 6228 -29637 6264
rect -32220 -1278 -32202 6228
rect -30789 5670 -30555 5688
rect -29871 5652 -29718 5670
rect -27882 5670 -27864 7767
rect -29007 5643 -28836 5670
rect -28332 5652 -27864 5670
rect -28656 5508 -28638 5535
rect -28656 5490 -28566 5508
rect -28584 5454 -28566 5490
rect -28584 5436 -28008 5454
rect -33309 -1305 -32202 -1278
rect -32130 4365 -29610 4383
rect -35307 -1557 -33705 -1539
rect -32130 -1809 -32112 4365
rect -30915 3807 -30834 3825
rect -30915 2610 -30897 3807
rect -30699 3735 -30555 3744
rect -29871 3717 -29718 3735
rect -27882 3735 -27864 5652
rect -29007 3708 -28836 3735
rect -28332 3717 -27864 3735
rect -28350 3708 -28332 3717
rect -28656 3573 -28638 3609
rect -28656 3555 -28566 3573
rect -28584 3492 -28566 3555
rect -28584 3474 -28260 3492
rect -28278 2610 -28260 3474
rect -30915 2592 -28260 2610
rect -33309 -1836 -32112 -1809
rect -31284 63 -30195 81
rect -35181 -2106 -33705 -2088
rect -34551 -2655 -33696 -2628
rect -34713 -3123 -33696 -3087
rect -33696 -3600 -33678 -3591
rect -34893 -3627 -33678 -3600
rect -33309 -3843 -31806 -3816
rect -33696 -4104 -33678 -4095
rect -35001 -4131 -33678 -4104
rect -31284 -4662 -31266 63
rect -30843 -4617 -30825 -108
rect -29943 -171 -29925 -27
rect -29403 -27 -29151 0
rect -29403 -171 -29385 -27
rect -29943 -189 -29385 -171
rect -29268 -837 -29160 -810
rect -30672 -882 -30195 -864
rect -29934 -1107 -29916 -972
rect -29268 -1107 -29250 -837
rect -29934 -1125 -29250 -1107
rect -26946 -1188 -26928 -810
rect -26856 -1593 -26838 -792
rect -29277 -1683 -29178 -1656
rect -29988 -2133 -29970 -2052
rect -29943 -2133 -29925 -2034
rect -29277 -2133 -29259 -1683
rect -29997 -2169 -29961 -2133
rect -29943 -2151 -29916 -2133
rect -29898 -2151 -29259 -2133
rect -29988 -2268 -29970 -2169
rect -28566 -2268 -28548 -1620
rect -29988 -2286 -28548 -2268
rect -29331 -2979 -29241 -2952
rect -29943 -3429 -29925 -3330
rect -29331 -3429 -29313 -2979
rect -29943 -3447 -29313 -3429
rect -29898 -3645 -29880 -3447
rect -30735 -3663 -29880 -3645
rect -29790 -3726 -29772 -3672
rect -30753 -3744 -29772 -3726
rect -29943 -4500 -29925 -4356
rect -29403 -4356 -29151 -4329
rect -29403 -4500 -29385 -4356
rect -29943 -4518 -29385 -4500
rect -29943 -4617 -29925 -4518
rect -30843 -4635 -29925 -4617
rect -31284 -4680 -30915 -4662
rect -31284 -6579 -31266 -4680
rect -30843 -5544 -30825 -4635
rect -29268 -5166 -29160 -5139
rect -29934 -5436 -29916 -5301
rect -29268 -5436 -29250 -5166
rect -29934 -5454 -29250 -5436
rect -29934 -5616 -29916 -5454
rect -26946 -5517 -26928 -5139
rect -30942 -5634 -29916 -5616
rect -26856 -5922 -26838 -5121
rect -29277 -6012 -29178 -5985
rect -30240 -6786 -30222 -6444
rect -29988 -6462 -29970 -6381
rect -29943 -6444 -29925 -6363
rect -29997 -6498 -29961 -6462
rect -29277 -6462 -29259 -6012
rect -29925 -6480 -29259 -6462
rect -29988 -6597 -29970 -6498
rect -28566 -6597 -28548 -5949
rect -29988 -6615 -28548 -6597
rect -31266 -6813 -30879 -6786
rect -30861 -6813 -30222 -6786
rect -29331 -7308 -29241 -7281
rect -29943 -7758 -29925 -7659
rect -29331 -7758 -29313 -7308
rect -29943 -7776 -29313 -7758
rect -29331 -8001 -29313 -7776
rect -31149 -8010 -29313 -8001
rect -31167 -8019 -29313 -8010
rect -35649 -8478 -34254 -8460
rect -35496 -8955 -34245 -8937
rect -34209 -8955 -33687 -8937
rect -35370 -9414 -34335 -9396
rect -34308 -9414 -33660 -9396
rect -35199 -9954 -34461 -9936
rect -34416 -9954 -33687 -9936
rect -34542 -10413 -33687 -10395
rect -34686 -10881 -33687 -10863
rect -34875 -11313 -33687 -11295
rect -31167 -11574 -31149 -8019
rect -30186 -9423 -30168 -9108
rect -30780 -9441 -30168 -9423
rect -30186 -10377 -30168 -10053
rect -30942 -10395 -30168 -10377
rect -36045 -11637 -35910 -11619
rect -36045 -12222 -36027 -11637
rect -35019 -11898 -33678 -11880
rect -36027 -12249 -35973 -12222
rect -35991 -12519 -35973 -12249
rect -31167 -12303 -31149 -11628
rect -31167 -12321 -30195 -12303
rect -35991 -12537 -35910 -12519
rect -31707 -14166 -31689 -14139
rect -32166 -14184 -31689 -14166
rect -32166 -14382 -32148 -14184
rect -33291 -14409 -32148 -14382
rect -32139 -14607 -31707 -14589
rect -32139 -14877 -32121 -14607
rect -33291 -14904 -32121 -14877
rect -32031 -15039 -31707 -15021
rect -32031 -15291 -32013 -15039
rect -33291 -15318 -32013 -15291
rect -31707 -15822 -31689 -15534
rect -33291 -15849 -31689 -15822
<< m123contact >>
rect -29538 10458 -29520 10494
rect -29538 9765 -29520 9801
rect -30348 9738 -30330 9765
rect -33696 -630 -33678 -594
rect -33705 -702 -33660 -675
rect -29538 8361 -29520 8388
rect -30348 7641 -30330 7677
rect -29538 7668 -29520 7704
rect -29538 6219 -29511 6291
rect -29538 5553 -29511 5589
rect -30348 5526 -30330 5553
rect -35397 -1557 -35361 -1539
rect -29538 4347 -29511 4383
rect -30348 3591 -30330 3627
rect -29538 3618 -29511 3654
rect -29376 288 -29358 315
rect -35298 -2115 -35262 -2079
rect -33354 -2403 -33309 -2376
rect -34650 -2655 -34605 -2628
rect -33345 -2898 -33309 -2871
rect -34794 -3123 -34776 -3087
rect -33345 -3312 -33309 -3285
rect -34974 -3627 -34956 -3600
rect -31698 -3861 -31680 -3771
rect -35163 -4131 -35127 -4104
rect -30636 -378 -30618 -333
rect -30465 -351 -30429 -333
rect -27882 -432 -27864 -387
rect -29385 -657 -29358 -630
rect -29412 -1674 -29385 -1647
rect -28404 -1647 -28377 -1620
rect -28143 -1647 -28116 -1620
rect -30816 -2340 -30789 -2322
rect -30726 -2412 -30708 -2385
rect -30483 -2403 -30429 -2385
rect -28701 -2943 -28674 -2916
rect -28557 -2943 -28530 -2916
rect -28431 -2943 -28404 -2916
rect -28296 -2943 -28269 -2916
rect -29988 -3348 -29970 -3321
rect -29790 -3627 -29772 -3609
rect -30816 -3663 -30789 -3645
rect -29376 -4041 -29358 -4014
rect -27882 -4761 -27864 -4716
rect -29385 -4986 -29358 -4959
rect -29412 -6003 -29385 -5976
rect -28404 -5976 -28377 -5949
rect -28143 -5976 -28116 -5949
rect -31437 -6813 -31419 -6786
rect -28701 -7272 -28674 -7245
rect -28557 -7272 -28530 -7245
rect -28431 -7272 -28404 -7245
rect -28296 -7272 -28269 -7245
rect -29988 -7677 -29970 -7650
rect -35676 -8424 -35658 -8361
rect -34164 -8478 -34110 -8460
rect -33687 -8487 -33651 -8451
rect -35523 -8919 -35496 -8883
rect -34236 -9027 -34218 -8973
rect -31437 -9117 -31419 -9036
rect -35397 -9369 -35361 -9324
rect -34335 -9450 -34308 -9423
rect -31284 -9486 -31266 -9468
rect -31374 -9711 -31356 -9648
rect -35289 -9963 -35271 -9927
rect -34461 -10044 -34425 -9990
rect -34641 -10422 -34614 -10386
rect -31230 -10431 -31212 -10413
rect -34794 -10890 -34776 -10854
rect -34983 -11322 -34947 -11286
rect -29781 -9486 -29763 -9468
rect -29781 -10431 -29763 -10413
rect -35748 -11655 -35712 -11637
rect -33975 -11745 -33957 -11709
rect -35154 -11907 -35127 -11871
rect -35757 -12123 -35703 -12105
rect -33336 -12474 -33291 -12447
rect -36063 -12573 -36009 -12546
rect -33975 -12645 -33957 -12591
rect -33687 -12681 -33642 -12645
rect -31374 -12663 -31356 -12618
rect -33336 -12969 -33291 -12942
rect -33678 -13158 -33660 -13140
rect -33327 -13383 -33291 -13356
rect -33687 -13662 -33642 -13617
rect -33336 -13914 -33291 -13887
rect -33687 -14139 -33651 -14112
rect -31869 -14157 -31851 -14139
rect -33678 -14643 -33660 -14607
rect -31869 -14634 -31851 -14616
rect -31869 -15003 -31851 -14976
rect -33678 -15120 -33660 -15093
rect -31869 -15516 -31851 -15480
rect -33687 -15570 -33651 -15525
rect -33678 -16092 -33660 -16056
<< metal3 >>
rect -29538 9801 -29520 10458
rect -30348 9027 -30330 9738
rect -32049 9009 -30330 9027
rect -35676 -621 -33696 -603
rect -35676 -8361 -35658 -621
rect -35523 -693 -33705 -675
rect -35523 -8883 -35505 -693
rect -35388 -9324 -35370 -1557
rect -35289 -9927 -35271 -2115
rect -32049 -2376 -32031 9009
rect -29538 7704 -29520 8361
rect -33309 -2403 -32031 -2376
rect -31959 6966 -31941 6975
rect -30348 6966 -30330 7641
rect -31959 6948 -30330 6966
rect -35748 -11817 -35730 -11655
rect -36027 -11835 -35730 -11817
rect -36027 -12204 -36009 -11835
rect -35154 -11871 -35136 -4131
rect -34974 -11286 -34956 -3627
rect -34794 -10854 -34776 -3123
rect -34632 -10386 -34614 -2655
rect -31959 -2871 -31941 6948
rect -29538 5589 -29511 6219
rect -29538 5526 -29511 5553
rect -30348 4788 -30330 5526
rect -33309 -2898 -31941 -2871
rect -31815 4770 -30330 4788
rect -31815 -3285 -31797 4770
rect -29538 3654 -29511 4347
rect -29538 3591 -29511 3618
rect -30348 3438 -30330 3591
rect -33309 -3312 -31797 -3285
rect -31698 3420 -30330 3438
rect -31698 -3771 -31680 3420
rect -30528 630 -29259 648
rect -31437 -2340 -30816 -2322
rect -31437 -6786 -31419 -2340
rect -34110 -8478 -33687 -8460
rect -35757 -12204 -35739 -12123
rect -36027 -12222 -35739 -12204
rect -36027 -12546 -36009 -12222
rect -35154 -16101 -35136 -11907
rect -34974 -15525 -34956 -11322
rect -34794 -15102 -34776 -10890
rect -34632 -14616 -34614 -10422
rect -34452 -14148 -34434 -10044
rect -34335 -13626 -34317 -9450
rect -34236 -13140 -34218 -9027
rect -34164 -12654 -34146 -8478
rect -31437 -9036 -31419 -6813
rect -31374 -3663 -30816 -3645
rect -31374 -7938 -31356 -3663
rect -30726 -6732 -30708 -2412
rect -30636 -5571 -30618 -378
rect -30528 -3690 -30510 630
rect -29376 270 -29358 288
rect -29277 270 -29259 630
rect -29376 252 -29259 270
rect -30429 -351 -29583 -333
rect -29601 -414 -29583 -351
rect -29376 -369 -29358 252
rect -29376 -387 -27864 -369
rect -29601 -432 -29268 -414
rect -29376 -684 -29358 -657
rect -29286 -684 -29268 -432
rect -29376 -702 -29268 -684
rect -29376 -1170 -29358 -702
rect -29376 -1188 -28422 -1170
rect -28440 -1620 -28422 -1188
rect -28116 -1341 -28098 -387
rect -28188 -1359 -28098 -1341
rect -28188 -1620 -28170 -1359
rect -28440 -1647 -28404 -1620
rect -28188 -1647 -28143 -1620
rect -29385 -1674 -29349 -1647
rect -29367 -2385 -29349 -1674
rect -30429 -2403 -29349 -2385
rect -29367 -2601 -29349 -2403
rect -28440 -2601 -28422 -1647
rect -29367 -2619 -28737 -2601
rect -28755 -2916 -28737 -2619
rect -28611 -2619 -28422 -2601
rect -28611 -2916 -28593 -2619
rect -28188 -2646 -28170 -1647
rect -28458 -2664 -28170 -2646
rect -28458 -2916 -28440 -2664
rect -28755 -2943 -28701 -2916
rect -28611 -2943 -28557 -2916
rect -28458 -2943 -28431 -2916
rect -28341 -2943 -28296 -2916
rect -29988 -3609 -29970 -3348
rect -28341 -3609 -28323 -2943
rect -29988 -3627 -29790 -3609
rect -29772 -3627 -28323 -3609
rect -30528 -3708 -29358 -3690
rect -29376 -4014 -29358 -3708
rect -29376 -4698 -29358 -4041
rect -29376 -4716 -27864 -4698
rect -29376 -5499 -29358 -4986
rect -29376 -5517 -28422 -5499
rect -29376 -5571 -29358 -5517
rect -30636 -5589 -29358 -5571
rect -28440 -5949 -28422 -5517
rect -28116 -5670 -28098 -4716
rect -28188 -5688 -28098 -5670
rect -28188 -5949 -28170 -5688
rect -28440 -5976 -28404 -5949
rect -28188 -5976 -28143 -5949
rect -29385 -6003 -29349 -5976
rect -29367 -6732 -29349 -6003
rect -30726 -6750 -29349 -6732
rect -29367 -6930 -29349 -6750
rect -28440 -6930 -28422 -5976
rect -29367 -6948 -28737 -6930
rect -28755 -7245 -28737 -6948
rect -28611 -6948 -28422 -6930
rect -28611 -7245 -28593 -6948
rect -28188 -6975 -28170 -5976
rect -28458 -6993 -28170 -6975
rect -28458 -7245 -28440 -6993
rect -28755 -7272 -28701 -7245
rect -28611 -7272 -28557 -7245
rect -28458 -7272 -28431 -7245
rect -28341 -7272 -28296 -7245
rect -29988 -7938 -29970 -7677
rect -28341 -7938 -28323 -7272
rect -31374 -7956 -31284 -7938
rect -31266 -7956 -28323 -7938
rect -31374 -9648 -31356 -7956
rect -31266 -9486 -29781 -9468
rect -33975 -12591 -33957 -11745
rect -33291 -12474 -32553 -12447
rect -34164 -12672 -33687 -12654
rect -33291 -12969 -32742 -12942
rect -34236 -13158 -33678 -13140
rect -33291 -13383 -32931 -13356
rect -34335 -13644 -33687 -13626
rect -33291 -13914 -33057 -13887
rect -33678 -14148 -33660 -14139
rect -34452 -14166 -33660 -14148
rect -34632 -14643 -33678 -14616
rect -34794 -15120 -33678 -15102
rect -34974 -15561 -33687 -15525
rect -33075 -15534 -33057 -13914
rect -32949 -15012 -32931 -13383
rect -32760 -14616 -32742 -12969
rect -32571 -14139 -32553 -12474
rect -31374 -12618 -31356 -9711
rect -31212 -10431 -29781 -10413
rect -32571 -14157 -31869 -14139
rect -32760 -14634 -31869 -14616
rect -31869 -15012 -31851 -15003
rect -32949 -15030 -31851 -15012
rect -31869 -15534 -31851 -15516
rect -33075 -15561 -31851 -15534
rect -33678 -16101 -33660 -16092
rect -35154 -16119 -33660 -16101
<< labels >>
rlabel polysilicon -36297 -12168 -36297 -12168 1 s0
rlabel polysilicon -36243 -12564 -36243 -12564 1 s1
rlabel metal1 -36198 -11772 -36198 -11772 1 vdd
rlabel polycontact -35298 -12906 -35298 -12906 1 D3
rlabel polycontact -35298 -12492 -35298 -12492 1 D2
rlabel polycontact -35316 -12051 -35316 -12051 1 D1
rlabel polycontact -35307 -11574 -35307 -11574 1 D0
rlabel metal1 -36081 -12240 -36081 -12240 1 s0_not
rlabel metal1 -36072 -12564 -36072 -12564 1 s1_not
rlabel polysilicon -33669 -12537 -33669 -12537 1 a3
rlabel polysilicon -33669 -13023 -33669 -13023 1 a2
rlabel polysilicon -33669 -13437 -33669 -13437 1 a1
rlabel polysilicon -33669 -13968 -33669 -13968 1 a0
rlabel m123contact -33318 -13905 -33318 -13905 1 and_a0
rlabel m123contact -33318 -13374 -33318 -13374 1 and_a1
rlabel m123contact -33318 -12960 -33318 -12960 1 and_a2
rlabel m123contact -33309 -12456 -33309 -12456 1 and_a3
rlabel polysilicon -33669 -14454 -33669 -14454 1 b3
rlabel polysilicon -33669 -14958 -33669 -14958 1 b2
rlabel polysilicon -33669 -15372 -33669 -15372 1 b1
rlabel polysilicon -33669 -15903 -33669 -15903 1 b0
rlabel m2contact -33318 -15840 -33318 -15840 1 and_b0
rlabel m2contact -33309 -15309 -33309 -15309 1 and_b1
rlabel m2contact -33300 -14895 -33300 -14895 1 and_b2
rlabel m2contact -33309 -14400 -33309 -14400 1 and_b3
rlabel polycontact -33309 -8244 -33309 -8244 1 comp_a3
rlabel polycontact -33309 -8730 -33309 -8730 1 comp_a2
rlabel polycontact -33309 -9144 -33309 -9144 1 comp_a1
rlabel polycontact -33309 -9684 -33309 -9684 1 comp_a0
rlabel polycontact -33318 -10161 -33318 -10161 1 comp_b3
rlabel polycontact -33309 -10656 -33309 -10656 1 comp_b2
rlabel polycontact -33309 -11061 -33309 -11061 1 comp_b1
rlabel polycontact -33309 -11601 -33309 -11601 1 comp_b0
rlabel metal1 -31347 -15246 -31347 -15246 1 and_oper_out0
rlabel metal1 -31347 -14778 -31347 -14778 1 and_oper_out1
rlabel metal1 -31338 -14391 -31338 -14391 1 and_oper_out2
rlabel metal1 -31338 -13914 -31338 -13914 1 and_oper_out3
rlabel metal1 -29394 -2952 -29394 -2952 1 x0
rlabel m123contact -29403 -1656 -29403 -1656 1 x1
rlabel metal1 -29394 -639 -29394 -639 1 x2
rlabel metal1 -29403 306 -29403 306 1 x3
rlabel metal1 -29052 -9 -29052 -9 1 a3_not
rlabel metal1 -28215 36 -28215 36 1 AlessB_3
rlabel metal1 -29070 -810 -29070 -810 1 a2_not
rlabel metal1 -27459 -774 -27459 -774 1 AlessB_2
rlabel metal1 -26649 -828 -26649 -828 7 AlessB
rlabel metal1 -29088 -1656 -29088 -1656 1 a1_not
rlabel metal1 -27801 -1602 -27801 -1602 1 AlessB_1
rlabel metal1 -29133 -2952 -29133 -2952 1 a0_not
rlabel metal1 -27945 -2898 -27945 -2898 1 AlessB_0
rlabel metal1 -29052 -4329 -29052 -4329 1 b3_not
rlabel metal1 -29070 -5139 -29070 -5139 1 b2_not
rlabel metal1 -29088 -5985 -29088 -5985 1 b1_not
rlabel metal1 -29133 -7290 -29133 -7290 1 b0_not
rlabel metal1 -27954 -7218 -27954 -7218 1 AmoreB_0
rlabel metal1 -27783 -5931 -27783 -5931 1 AmoreB_1
rlabel metal1 -27450 -5103 -27450 -5103 1 AmoreB_2
rlabel metal1 -28206 -4302 -28206 -4302 1 AmoreB_3
rlabel metal1 -26640 -5157 -26640 -5157 7 AmoreB
rlabel metal1 -28269 -5967 -28269 -5967 1 temp_more
rlabel metal1 -28269 -1638 -28269 -1638 1 temp_less
rlabel polycontact -27297 -9882 -27297 -9882 1 k
rlabel polysilicon -27630 -9918 -27630 -9918 1 temp
rlabel metal1 -26307 -9828 -26307 -9828 1 AequalsB
rlabel polysilicon -26658 -9900 -26658 -9900 1 equals_d
rlabel polysilicon -34074 -1170 -34074 -1170 1 D
rlabel m2contact -33336 -378 -33336 -378 1 adsub_a3
rlabel m2contact -33327 -882 -33327 -882 1 adsub_a2
rlabel m2contact -33327 -1296 -33327 -1296 1 adsub_a1
rlabel m123contact -33327 -2394 -33327 -2394 1 adsub_b3
rlabel m123contact -33327 -2880 -33327 -2880 1 adsub_b2
rlabel m123contact -33336 -3294 -33336 -3294 1 adsub_b1
rlabel m2contact -33327 -3825 -33327 -3825 1 adsub_b0
rlabel polysilicon -28296 4032 -28296 4032 7 sum0
rlabel metal1 -29376 2736 -29376 2736 1 carry0
rlabel polysilicon -28287 5967 -28287 5967 1 sum1
rlabel polycontact -29385 4671 -29385 4671 1 carry1
rlabel polysilicon -28305 8082 -28305 8082 1 sum2
rlabel metal1 -29385 6786 -29385 6786 1 carry2
rlabel polysilicon -28296 10179 -28296 10179 1 sum3
rlabel metal1 -29385 8883 -29385 8883 1 carry3
rlabel metal1 -36189 -12888 -36189 -12888 1 gnd!
rlabel m2contact -33327 -1827 -33327 -1827 1 adsub_a0
<< end >>
