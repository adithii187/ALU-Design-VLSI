magic
tech scmos
magscale 9 1
timestamp 1700400098
<< nwell >>
rect 17 -26 56 -13
<< ntransistor >>
rect 24 -37 26 -34
rect 34 -37 36 -34
rect 48 -37 50 -34
<< ptransistor >>
rect 24 -24 26 -19
rect 34 -24 36 -19
rect 48 -24 50 -19
<< ndiffusion >>
rect 20 -36 21 -34
rect 23 -36 24 -34
rect 20 -37 24 -36
rect 26 -36 27 -34
rect 26 -37 29 -36
rect 30 -36 31 -34
rect 33 -36 34 -34
rect 30 -37 34 -36
rect 36 -36 37 -34
rect 36 -37 39 -36
rect 44 -36 45 -34
rect 47 -36 48 -34
rect 44 -37 48 -36
rect 50 -36 51 -34
rect 53 -36 54 -34
rect 50 -37 54 -36
<< pdiffusion >>
rect 19 -20 24 -19
rect 19 -22 20 -20
rect 22 -22 24 -20
rect 19 -24 24 -22
rect 26 -24 34 -19
rect 36 -21 39 -19
rect 36 -23 37 -21
rect 36 -24 39 -23
rect 44 -20 48 -19
rect 44 -22 45 -20
rect 47 -22 48 -20
rect 44 -24 48 -22
rect 50 -21 54 -19
rect 50 -23 51 -21
rect 53 -23 54 -21
rect 50 -24 54 -23
<< ndcontact >>
rect 21 -36 23 -34
rect 27 -36 29 -34
rect 31 -36 33 -34
rect 37 -36 39 -34
rect 45 -36 47 -34
rect 51 -36 53 -34
<< pdcontact >>
rect 20 -22 22 -20
rect 37 -23 39 -21
rect 45 -22 47 -20
rect 51 -23 53 -21
<< polysilicon >>
rect 24 -19 26 -17
rect 34 -19 36 -17
rect 48 -19 50 -17
rect 24 -34 26 -24
rect 34 -34 36 -24
rect 48 -29 50 -24
rect 49 -31 50 -29
rect 48 -34 50 -31
rect 24 -38 26 -37
rect 34 -38 36 -37
rect 48 -38 50 -37
<< polycontact >>
rect 48 -31 49 -29
<< metal1 >>
rect 20 -16 50 -14
rect 20 -20 22 -16
rect 45 -20 47 -16
rect 37 -29 39 -23
rect 51 -29 53 -23
rect 27 -31 48 -29
rect 51 -31 56 -29
rect 27 -34 29 -31
rect 37 -34 39 -31
rect 51 -34 53 -31
rect 21 -39 23 -36
rect 31 -39 33 -36
rect 45 -39 47 -36
rect 19 -41 47 -39
<< labels >>
rlabel metal1 31 -40 31 -40 1 gnd
rlabel metal1 34 -15 34 -15 5 vdd
rlabel metal1 54 -30 54 -30 7 out
rlabel polysilicon 25 -29 25 -29 1 a
rlabel polysilicon 35 -28 35 -28 1 b
<< end >>
