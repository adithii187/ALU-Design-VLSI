magic
tech scmos
magscale 9 1
timestamp 1700922776
<< nwell >>
rect -249 350 -237 425
rect -210 417 -189 422
rect -209 405 -192 417
rect -209 404 -202 405
rect -200 404 -192 405
rect -169 383 -148 388
rect -75 387 -54 393
rect -168 371 -151 383
rect -168 370 -161 371
rect -159 370 -151 371
rect -127 370 -91 380
rect -75 375 -58 387
rect -75 374 -68 375
rect -66 374 -58 375
rect -249 245 -237 320
rect -210 312 -189 317
rect -209 300 -192 312
rect -209 299 -202 300
rect -200 299 -192 300
rect -171 295 -150 298
rect -172 293 -150 295
rect -83 297 -62 303
rect 9 300 30 303
rect 9 298 61 300
rect 9 297 30 298
rect -170 281 -153 293
rect -170 280 -163 281
rect -161 280 -153 281
rect -135 280 -99 290
rect -83 285 -66 297
rect -83 284 -76 285
rect -74 284 -66 285
rect -43 280 -7 290
rect 9 285 26 297
rect 59 293 61 298
rect 9 284 16 285
rect 18 284 26 285
rect 57 280 115 293
rect 91 278 95 280
rect -119 209 -9 212
rect -249 132 -237 207
rect -120 206 -9 209
rect -210 199 -190 204
rect -173 199 -152 204
rect -209 187 -192 199
rect -209 186 -202 187
rect -200 186 -192 187
rect -172 187 -155 199
rect -119 194 -9 206
rect -172 186 -165 187
rect -163 186 -155 187
rect -136 65 -26 68
rect -249 -12 -237 63
rect -137 62 -26 65
rect -210 55 -190 60
rect -179 55 -158 60
rect -209 43 -192 55
rect -209 42 -202 43
rect -200 42 -192 43
rect -178 43 -161 55
rect -136 50 -26 62
rect -178 42 -171 43
rect -169 42 -161 43
<< ntransistor >>
rect -274 416 -268 418
rect -274 397 -268 399
rect -202 395 -200 398
rect -274 375 -268 377
rect -274 357 -268 359
rect -161 361 -159 364
rect -68 365 -66 368
rect -119 359 -117 362
rect -107 359 -106 362
rect -101 359 -99 362
rect -274 311 -268 313
rect -274 292 -268 294
rect -202 290 -200 293
rect -274 270 -268 272
rect -163 271 -161 274
rect -76 275 -74 278
rect 16 275 18 278
rect -127 269 -125 272
rect -115 269 -114 272
rect -109 269 -107 272
rect -35 269 -33 272
rect -17 269 -15 272
rect 63 269 65 272
rect 73 269 75 272
rect 83 269 85 272
rect 93 269 95 272
rect 107 269 109 272
rect -274 252 -268 254
rect -274 198 -268 200
rect -274 179 -268 181
rect -202 177 -200 180
rect -165 177 -163 180
rect -109 179 -107 182
rect -95 179 -93 182
rect -79 179 -77 182
rect -65 179 -63 182
rect -50 179 -48 182
rect -21 179 -19 182
rect -274 157 -268 159
rect -274 139 -268 141
rect -274 54 -268 56
rect -274 35 -268 37
rect -202 33 -200 36
rect -171 33 -169 36
rect -126 35 -124 38
rect -112 35 -110 38
rect -96 35 -94 38
rect -82 35 -80 38
rect -67 35 -65 38
rect -38 35 -36 38
rect -274 13 -268 15
rect -274 -5 -268 -3
<< ptransistor >>
rect -246 416 -239 418
rect -202 406 -200 412
rect -246 397 -239 399
rect -246 375 -239 377
rect -246 357 -239 359
rect -161 372 -159 378
rect -119 373 -117 378
rect -101 373 -99 378
rect -68 376 -66 382
rect -246 311 -239 313
rect -202 301 -200 307
rect -246 292 -239 294
rect -246 270 -239 272
rect -163 282 -161 288
rect -127 283 -125 288
rect -109 283 -107 288
rect -76 286 -74 292
rect -35 283 -33 288
rect -17 283 -15 288
rect 16 286 18 292
rect 63 282 65 287
rect 69 282 71 287
rect 73 282 75 287
rect 83 282 85 287
rect 93 282 95 287
rect 107 282 109 287
rect -246 252 -239 254
rect -246 198 -239 200
rect -109 196 -107 202
rect -95 196 -93 202
rect -79 196 -77 202
rect -65 196 -63 202
rect -50 196 -48 202
rect -21 196 -19 202
rect -202 188 -200 194
rect -165 188 -163 194
rect -246 179 -239 181
rect -246 157 -239 159
rect -246 139 -239 141
rect -246 54 -239 56
rect -126 52 -124 58
rect -112 52 -110 58
rect -96 52 -94 58
rect -82 52 -80 58
rect -67 52 -65 58
rect -38 52 -36 58
rect -202 44 -200 50
rect -171 44 -169 50
rect -246 35 -239 37
rect -246 13 -239 15
rect -246 -5 -239 -3
<< ndiffusion >>
rect -274 423 -268 424
rect -274 419 -273 423
rect -269 419 -268 423
rect -274 418 -268 419
rect -274 415 -268 416
rect -274 411 -273 415
rect -269 411 -268 415
rect -274 410 -268 411
rect -274 404 -268 405
rect -274 400 -273 404
rect -269 400 -268 404
rect -274 399 -268 400
rect -207 397 -202 398
rect -274 396 -268 397
rect -274 392 -273 396
rect -269 392 -268 396
rect -274 391 -268 392
rect -207 395 -206 397
rect -203 395 -202 397
rect -200 395 -198 398
rect -195 395 -194 398
rect -274 383 -268 384
rect -274 379 -273 383
rect -269 379 -268 383
rect -274 377 -268 379
rect -274 374 -268 375
rect -274 370 -273 374
rect -269 370 -268 374
rect -274 369 -268 370
rect -274 365 -268 366
rect -274 361 -273 365
rect -269 361 -268 365
rect -274 359 -268 361
rect -274 356 -268 357
rect -274 352 -273 356
rect -269 352 -268 356
rect -274 351 -268 352
rect -166 363 -161 364
rect -166 361 -165 363
rect -162 361 -161 363
rect -159 361 -157 364
rect -154 361 -153 364
rect -73 367 -68 368
rect -73 365 -72 367
rect -69 365 -68 367
rect -66 365 -64 368
rect -61 365 -60 368
rect -123 361 -119 362
rect -123 359 -122 361
rect -120 359 -119 361
rect -117 359 -107 362
rect -106 359 -101 362
rect -99 360 -98 362
rect -96 360 -95 362
rect -99 359 -95 360
rect -274 318 -268 319
rect -274 314 -273 318
rect -269 314 -268 318
rect -274 313 -268 314
rect -274 310 -268 311
rect -274 306 -273 310
rect -269 306 -268 310
rect -274 305 -268 306
rect -274 299 -268 300
rect -274 295 -273 299
rect -269 295 -268 299
rect -274 294 -268 295
rect -207 292 -202 293
rect -274 291 -268 292
rect -274 287 -273 291
rect -269 287 -268 291
rect -274 286 -268 287
rect -207 290 -206 292
rect -203 290 -202 292
rect -200 290 -198 293
rect -195 290 -194 293
rect -274 278 -268 279
rect -274 274 -273 278
rect -269 274 -268 278
rect -274 272 -268 274
rect -274 269 -268 270
rect -274 265 -273 269
rect -269 265 -268 269
rect -274 264 -268 265
rect -168 273 -163 274
rect -168 271 -167 273
rect -164 271 -163 273
rect -161 271 -159 274
rect -156 271 -155 274
rect -81 277 -76 278
rect -81 275 -80 277
rect -77 275 -76 277
rect -74 275 -72 278
rect -69 275 -68 278
rect 11 277 16 278
rect 11 275 12 277
rect 15 275 16 277
rect 18 275 20 278
rect 23 275 24 278
rect -131 271 -127 272
rect -131 269 -130 271
rect -128 269 -127 271
rect -125 269 -115 272
rect -114 269 -109 272
rect -107 270 -106 272
rect -104 270 -103 272
rect -107 269 -103 270
rect -39 271 -35 272
rect -39 269 -38 271
rect -36 269 -35 271
rect -33 269 -17 272
rect -15 270 -14 272
rect -12 270 -11 272
rect -15 269 -11 270
rect 58 270 59 272
rect 61 270 63 272
rect 58 269 63 270
rect 65 270 66 272
rect 65 269 68 270
rect 69 270 70 272
rect 72 270 73 272
rect 69 269 73 270
rect 75 270 76 272
rect 75 269 78 270
rect 79 270 80 272
rect 82 270 83 272
rect 79 269 83 270
rect 85 270 86 272
rect 85 269 88 270
rect 89 270 90 272
rect 92 270 93 272
rect 89 269 93 270
rect 95 270 96 272
rect 95 269 98 270
rect 103 270 104 272
rect 106 270 107 272
rect 103 269 107 270
rect 109 270 110 272
rect 112 270 113 272
rect 109 269 113 270
rect -274 260 -268 261
rect -274 256 -273 260
rect -269 256 -268 260
rect -274 254 -268 256
rect -274 251 -268 252
rect -274 247 -273 251
rect -269 247 -268 251
rect -274 246 -268 247
rect -274 205 -268 206
rect -274 201 -273 205
rect -269 201 -268 205
rect -274 200 -268 201
rect -274 197 -268 198
rect -274 193 -273 197
rect -269 193 -268 197
rect -274 192 -268 193
rect -274 186 -268 187
rect -274 182 -273 186
rect -269 182 -268 186
rect -274 181 -268 182
rect -207 179 -202 180
rect -274 178 -268 179
rect -274 174 -273 178
rect -269 174 -268 178
rect -274 173 -268 174
rect -207 177 -206 179
rect -203 177 -202 179
rect -200 177 -198 180
rect -195 177 -194 180
rect -170 179 -165 180
rect -170 177 -169 179
rect -166 177 -165 179
rect -163 177 -161 180
rect -158 177 -157 180
rect -114 179 -113 182
rect -110 179 -109 182
rect -107 179 -95 182
rect -93 179 -79 182
rect -77 179 -65 182
rect -63 179 -50 182
rect -48 179 -44 182
rect -41 179 -33 182
rect -27 179 -25 182
rect -22 179 -21 182
rect -19 179 -18 182
rect -15 179 -14 182
rect -274 165 -268 166
rect -274 161 -273 165
rect -269 161 -268 165
rect -274 159 -268 161
rect -274 156 -268 157
rect -274 152 -273 156
rect -269 152 -268 156
rect -274 151 -268 152
rect -274 147 -268 148
rect -274 143 -273 147
rect -269 143 -268 147
rect -274 141 -268 143
rect -274 138 -268 139
rect -274 134 -273 138
rect -269 134 -268 138
rect -274 133 -268 134
rect -274 61 -268 62
rect -274 57 -273 61
rect -269 57 -268 61
rect -274 56 -268 57
rect -274 53 -268 54
rect -274 49 -273 53
rect -269 49 -268 53
rect -274 48 -268 49
rect -274 42 -268 43
rect -274 38 -273 42
rect -269 38 -268 42
rect -274 37 -268 38
rect -207 35 -202 36
rect -274 34 -268 35
rect -274 30 -273 34
rect -269 30 -268 34
rect -274 29 -268 30
rect -207 33 -206 35
rect -203 33 -202 35
rect -200 33 -198 36
rect -195 33 -194 36
rect -176 35 -171 36
rect -176 33 -175 35
rect -172 33 -171 35
rect -169 33 -167 36
rect -164 33 -163 36
rect -131 35 -130 38
rect -127 35 -126 38
rect -124 35 -112 38
rect -110 35 -96 38
rect -94 35 -82 38
rect -80 35 -67 38
rect -65 35 -61 38
rect -58 35 -50 38
rect -44 35 -42 38
rect -39 35 -38 38
rect -36 35 -35 38
rect -32 35 -31 38
rect -274 21 -268 22
rect -274 17 -273 21
rect -269 17 -268 21
rect -274 15 -268 17
rect -274 12 -268 13
rect -274 8 -273 12
rect -269 8 -268 12
rect -274 7 -268 8
rect -274 3 -268 4
rect -274 -1 -273 3
rect -269 -1 -268 3
rect -274 -3 -268 -1
rect -274 -6 -268 -5
rect -274 -10 -273 -6
rect -269 -10 -268 -6
rect -274 -11 -268 -10
<< pdiffusion >>
rect -246 423 -239 424
rect -246 419 -245 423
rect -241 419 -239 423
rect -246 418 -239 419
rect -246 415 -239 416
rect -246 411 -245 415
rect -241 411 -239 415
rect -246 410 -239 411
rect -246 404 -239 405
rect -246 400 -245 404
rect -241 400 -239 404
rect -246 399 -239 400
rect -207 409 -206 412
rect -203 409 -202 412
rect -207 406 -202 409
rect -200 411 -194 412
rect -200 408 -198 411
rect -195 408 -194 411
rect -200 406 -194 408
rect -246 396 -239 397
rect -246 392 -245 396
rect -241 392 -239 396
rect -246 391 -239 392
rect -246 383 -239 384
rect -246 379 -245 383
rect -241 379 -239 383
rect -246 377 -239 379
rect -246 374 -239 375
rect -246 370 -245 374
rect -241 370 -239 374
rect -246 369 -239 370
rect -246 365 -239 366
rect -246 361 -245 365
rect -241 361 -239 365
rect -246 359 -239 361
rect -246 356 -239 357
rect -246 352 -245 356
rect -241 352 -239 356
rect -246 351 -239 352
rect -73 379 -72 382
rect -69 379 -68 382
rect -166 375 -165 378
rect -162 375 -161 378
rect -166 372 -161 375
rect -159 377 -153 378
rect -159 374 -157 377
rect -154 374 -153 377
rect -159 372 -153 374
rect -123 377 -119 378
rect -123 375 -122 377
rect -120 375 -119 377
rect -123 373 -119 375
rect -117 376 -110 378
rect -117 374 -116 376
rect -114 374 -110 376
rect -117 373 -110 374
rect -106 377 -101 378
rect -106 375 -105 377
rect -103 375 -101 377
rect -106 373 -101 375
rect -99 377 -95 378
rect -99 375 -98 377
rect -96 375 -95 377
rect -73 376 -68 379
rect -66 381 -60 382
rect -66 378 -64 381
rect -61 378 -60 381
rect -66 376 -60 378
rect -99 373 -95 375
rect -246 318 -239 319
rect -246 314 -245 318
rect -241 314 -239 318
rect -246 313 -239 314
rect -246 310 -239 311
rect -246 306 -245 310
rect -241 306 -239 310
rect -246 305 -239 306
rect -246 299 -239 300
rect -246 295 -245 299
rect -241 295 -239 299
rect -246 294 -239 295
rect -207 304 -206 307
rect -203 304 -202 307
rect -207 301 -202 304
rect -200 306 -194 307
rect -200 303 -198 306
rect -195 303 -194 306
rect -200 301 -194 303
rect -246 291 -239 292
rect -246 287 -245 291
rect -241 287 -239 291
rect -81 289 -80 292
rect -77 289 -76 292
rect -246 286 -239 287
rect -246 278 -239 279
rect -246 274 -245 278
rect -241 274 -239 278
rect -246 272 -239 274
rect -246 269 -239 270
rect -246 265 -245 269
rect -241 265 -239 269
rect -168 285 -167 288
rect -164 285 -163 288
rect -168 282 -163 285
rect -161 287 -155 288
rect -161 284 -159 287
rect -156 284 -155 287
rect -161 282 -155 284
rect -131 287 -127 288
rect -131 285 -130 287
rect -128 285 -127 287
rect -131 283 -127 285
rect -125 286 -118 288
rect -125 284 -124 286
rect -122 284 -118 286
rect -125 283 -118 284
rect -114 287 -109 288
rect -114 285 -113 287
rect -111 285 -109 287
rect -114 283 -109 285
rect -107 287 -103 288
rect -107 285 -106 287
rect -104 285 -103 287
rect -81 286 -76 289
rect -74 291 -68 292
rect -74 288 -72 291
rect -69 288 -68 291
rect -74 286 -68 288
rect -39 287 -35 288
rect -107 283 -103 285
rect -39 285 -38 287
rect -36 285 -35 287
rect -39 283 -35 285
rect -33 286 -26 288
rect -33 284 -32 286
rect -30 284 -26 286
rect -33 283 -26 284
rect 11 289 12 292
rect 15 289 16 292
rect -22 287 -17 288
rect -22 285 -21 287
rect -19 285 -17 287
rect -22 283 -17 285
rect -15 287 -11 288
rect -15 285 -14 287
rect -12 285 -11 287
rect 11 286 16 289
rect 18 291 24 292
rect 18 288 20 291
rect 23 288 24 291
rect 18 286 24 288
rect 58 286 63 287
rect -15 283 -11 285
rect 58 284 59 286
rect 61 284 63 286
rect 58 282 63 284
rect 65 282 69 287
rect 71 282 73 287
rect 75 282 83 287
rect 85 282 93 287
rect 95 285 98 287
rect 95 283 96 285
rect 95 282 98 283
rect 103 286 107 287
rect 103 284 104 286
rect 106 284 107 286
rect 103 282 107 284
rect 109 285 113 287
rect 109 283 110 285
rect 112 283 113 285
rect 109 282 113 283
rect -246 264 -239 265
rect -246 260 -239 261
rect -246 256 -245 260
rect -241 256 -239 260
rect -246 254 -239 256
rect -246 251 -239 252
rect -246 247 -245 251
rect -241 247 -239 251
rect -246 246 -239 247
rect -246 205 -239 206
rect -246 201 -245 205
rect -241 201 -239 205
rect -246 200 -239 201
rect -246 197 -239 198
rect -246 193 -245 197
rect -241 193 -239 197
rect -246 192 -239 193
rect -246 186 -239 187
rect -246 182 -245 186
rect -241 182 -239 186
rect -246 181 -239 182
rect -114 201 -109 202
rect -114 198 -113 201
rect -110 198 -109 201
rect -114 196 -109 198
rect -107 200 -102 202
rect -107 197 -106 200
rect -103 197 -102 200
rect -107 196 -102 197
rect -100 201 -95 202
rect -100 198 -99 201
rect -96 198 -95 201
rect -100 196 -95 198
rect -93 200 -87 202
rect -93 197 -92 200
rect -89 197 -87 200
rect -93 196 -87 197
rect -85 201 -79 202
rect -85 198 -83 201
rect -80 198 -79 201
rect -85 196 -79 198
rect -77 200 -72 202
rect -77 197 -76 200
rect -73 197 -72 200
rect -77 196 -72 197
rect -70 201 -65 202
rect -70 198 -69 201
rect -66 198 -65 201
rect -70 196 -65 198
rect -63 200 -58 202
rect -63 197 -62 200
rect -59 197 -58 200
rect -63 196 -58 197
rect -56 201 -50 202
rect -56 198 -55 201
rect -52 198 -50 201
rect -56 196 -50 198
rect -48 200 -33 202
rect -48 197 -47 200
rect -44 197 -33 200
rect -48 196 -33 197
rect -27 199 -25 202
rect -22 199 -21 202
rect -27 196 -21 199
rect -19 200 -14 202
rect -19 197 -18 200
rect -15 197 -14 200
rect -19 196 -14 197
rect -207 191 -206 194
rect -203 191 -202 194
rect -207 188 -202 191
rect -200 193 -194 194
rect -200 190 -198 193
rect -195 190 -194 193
rect -200 188 -194 190
rect -170 191 -169 194
rect -166 191 -165 194
rect -170 188 -165 191
rect -163 193 -157 194
rect -163 190 -161 193
rect -158 190 -157 193
rect -163 188 -157 190
rect -246 178 -239 179
rect -246 174 -245 178
rect -241 174 -239 178
rect -246 173 -239 174
rect -246 165 -239 166
rect -246 161 -245 165
rect -241 161 -239 165
rect -246 159 -239 161
rect -246 156 -239 157
rect -246 152 -245 156
rect -241 152 -239 156
rect -246 151 -239 152
rect -246 147 -239 148
rect -246 143 -245 147
rect -241 143 -239 147
rect -246 141 -239 143
rect -246 138 -239 139
rect -246 134 -245 138
rect -241 134 -239 138
rect -246 133 -239 134
rect -246 61 -239 62
rect -246 57 -245 61
rect -241 57 -239 61
rect -246 56 -239 57
rect -246 53 -239 54
rect -246 49 -245 53
rect -241 49 -239 53
rect -246 48 -239 49
rect -246 42 -239 43
rect -246 38 -245 42
rect -241 38 -239 42
rect -246 37 -239 38
rect -131 57 -126 58
rect -131 54 -130 57
rect -127 54 -126 57
rect -131 52 -126 54
rect -124 56 -119 58
rect -124 53 -123 56
rect -120 53 -119 56
rect -124 52 -119 53
rect -117 57 -112 58
rect -117 54 -116 57
rect -113 54 -112 57
rect -117 52 -112 54
rect -110 56 -104 58
rect -110 53 -109 56
rect -106 53 -104 56
rect -110 52 -104 53
rect -102 57 -96 58
rect -102 54 -100 57
rect -97 54 -96 57
rect -102 52 -96 54
rect -94 56 -89 58
rect -94 53 -93 56
rect -90 53 -89 56
rect -94 52 -89 53
rect -87 57 -82 58
rect -87 54 -86 57
rect -83 54 -82 57
rect -87 52 -82 54
rect -80 56 -75 58
rect -80 53 -79 56
rect -76 53 -75 56
rect -80 52 -75 53
rect -73 57 -67 58
rect -73 54 -72 57
rect -69 54 -67 57
rect -73 52 -67 54
rect -65 56 -50 58
rect -65 53 -64 56
rect -61 53 -50 56
rect -65 52 -50 53
rect -44 55 -42 58
rect -39 55 -38 58
rect -44 52 -38 55
rect -36 56 -31 58
rect -36 53 -35 56
rect -32 53 -31 56
rect -36 52 -31 53
rect -207 47 -206 50
rect -203 47 -202 50
rect -207 44 -202 47
rect -200 49 -194 50
rect -200 46 -198 49
rect -195 46 -194 49
rect -200 44 -194 46
rect -176 47 -175 50
rect -172 47 -171 50
rect -176 44 -171 47
rect -169 49 -163 50
rect -169 46 -167 49
rect -164 46 -163 49
rect -169 44 -163 46
rect -246 34 -239 35
rect -246 30 -245 34
rect -241 30 -239 34
rect -246 29 -239 30
rect -246 21 -239 22
rect -246 17 -245 21
rect -241 17 -239 21
rect -246 15 -239 17
rect -246 12 -239 13
rect -246 8 -245 12
rect -241 8 -239 12
rect -246 7 -239 8
rect -246 3 -239 4
rect -246 -1 -245 3
rect -241 -1 -239 3
rect -246 -3 -239 -1
rect -246 -6 -239 -5
rect -246 -10 -245 -6
rect -241 -10 -239 -6
rect -246 -11 -239 -10
<< ndcontact >>
rect -273 419 -269 423
rect -273 411 -269 415
rect -273 400 -269 404
rect -273 392 -269 396
rect -206 394 -203 397
rect -198 395 -195 398
rect -273 379 -269 383
rect -273 370 -269 374
rect -273 361 -269 365
rect -273 352 -269 356
rect -165 360 -162 363
rect -157 361 -154 364
rect -72 364 -69 367
rect -64 365 -61 368
rect -122 359 -120 361
rect -98 360 -96 362
rect -273 314 -269 318
rect -273 306 -269 310
rect -273 295 -269 299
rect -273 287 -269 291
rect -206 289 -203 292
rect -198 290 -195 293
rect -273 274 -269 278
rect -273 265 -269 269
rect -167 270 -164 273
rect -159 271 -156 274
rect -80 274 -77 277
rect -72 275 -69 278
rect 12 274 15 277
rect 20 275 23 278
rect -130 269 -128 271
rect -106 270 -104 272
rect -38 269 -36 271
rect -14 270 -12 272
rect 59 270 61 272
rect 66 270 68 272
rect 70 270 72 272
rect 76 270 78 272
rect 80 270 82 272
rect 86 270 88 272
rect 90 270 92 272
rect 96 270 98 272
rect 104 270 106 272
rect 110 270 112 272
rect -273 256 -269 260
rect -273 247 -269 251
rect -273 201 -269 205
rect -273 193 -269 197
rect -273 182 -269 186
rect -273 174 -269 178
rect -206 176 -203 179
rect -198 177 -195 180
rect -169 176 -166 179
rect -161 177 -158 180
rect -113 179 -110 182
rect -44 179 -41 182
rect -25 179 -22 182
rect -18 179 -15 182
rect -273 161 -269 165
rect -273 152 -269 156
rect -273 143 -269 147
rect -273 134 -269 138
rect -273 57 -269 61
rect -273 49 -269 53
rect -273 38 -269 42
rect -273 30 -269 34
rect -206 32 -203 35
rect -198 33 -195 36
rect -175 32 -172 35
rect -167 33 -164 36
rect -130 35 -127 38
rect -61 35 -58 38
rect -42 35 -39 38
rect -35 35 -32 38
rect -273 17 -269 21
rect -273 8 -269 12
rect -273 -1 -269 3
rect -273 -10 -269 -6
<< pdcontact >>
rect -245 419 -241 423
rect -245 411 -241 415
rect -245 400 -241 404
rect -206 409 -203 412
rect -198 408 -195 411
rect -245 392 -241 396
rect -245 379 -241 383
rect -245 370 -241 374
rect -245 361 -241 365
rect -245 352 -241 356
rect -72 379 -69 382
rect -165 375 -162 378
rect -157 374 -154 377
rect -122 375 -120 377
rect -116 374 -114 376
rect -105 375 -103 377
rect -98 375 -96 377
rect -64 378 -61 381
rect -245 314 -241 318
rect -245 306 -241 310
rect -245 295 -241 299
rect -206 304 -203 307
rect -198 303 -195 306
rect -245 287 -241 291
rect -80 289 -77 292
rect -245 274 -241 278
rect -245 265 -241 269
rect -167 285 -164 288
rect -159 284 -156 287
rect -130 285 -128 287
rect -124 284 -122 286
rect -113 285 -111 287
rect -106 285 -104 287
rect -72 288 -69 291
rect -38 285 -36 287
rect -32 284 -30 286
rect 12 289 15 292
rect -21 285 -19 287
rect -14 285 -12 287
rect 20 288 23 291
rect 59 284 61 286
rect 96 283 98 285
rect 104 284 106 286
rect 110 283 112 285
rect -245 256 -241 260
rect -245 247 -241 251
rect -245 201 -241 205
rect -245 193 -241 197
rect -245 182 -241 186
rect -113 198 -110 201
rect -106 197 -103 200
rect -99 198 -96 201
rect -92 197 -89 200
rect -83 198 -80 201
rect -76 197 -73 200
rect -69 198 -66 201
rect -62 197 -59 200
rect -55 198 -52 201
rect -47 197 -44 200
rect -25 199 -22 202
rect -18 197 -15 200
rect -206 191 -203 194
rect -198 190 -195 193
rect -169 191 -166 194
rect -161 190 -158 193
rect -245 174 -241 178
rect -245 161 -241 165
rect -245 152 -241 156
rect -245 143 -241 147
rect -245 134 -241 138
rect -245 57 -241 61
rect -245 49 -241 53
rect -245 38 -241 42
rect -130 54 -127 57
rect -123 53 -120 56
rect -116 54 -113 57
rect -109 53 -106 56
rect -100 54 -97 57
rect -93 53 -90 56
rect -86 54 -83 57
rect -79 53 -76 56
rect -72 54 -69 57
rect -64 53 -61 56
rect -42 55 -39 58
rect -35 53 -32 56
rect -206 47 -203 50
rect -198 46 -195 49
rect -175 47 -172 50
rect -167 46 -164 49
rect -245 30 -241 34
rect -245 17 -241 21
rect -245 8 -241 12
rect -245 -1 -241 3
rect -245 -10 -241 -6
<< psubstratepcontact >>
rect -287 375 -283 379
rect -287 365 -283 369
rect -287 270 -283 274
rect -287 260 -283 264
rect -287 157 -283 161
rect -287 147 -283 151
rect -287 13 -283 17
rect -287 3 -283 7
<< nsubstratencontact >>
rect -232 375 -228 379
rect -232 365 -228 369
rect -232 270 -228 274
rect -232 260 -228 264
rect -232 157 -228 161
rect -232 147 -228 151
rect -232 13 -228 17
rect -232 3 -228 7
<< polysilicon >>
rect -280 428 -231 430
rect -280 418 -278 428
rect -297 416 -274 418
rect -268 416 -267 418
rect -265 416 -246 418
rect -239 416 -236 418
rect -297 345 -295 416
rect -265 399 -263 416
rect -233 399 -231 428
rect -202 412 -200 414
rect -202 402 -200 406
rect -292 397 -274 399
rect -268 397 -263 399
rect -250 397 -246 399
rect -239 397 -231 399
rect -226 399 -206 402
rect -201 399 -200 402
rect -202 398 -200 399
rect -292 359 -290 397
rect -202 393 -200 395
rect -260 377 -256 380
rect -281 375 -274 377
rect -268 375 -246 377
rect -239 375 -234 377
rect -259 367 -257 375
rect -260 359 -256 364
rect -292 357 -274 359
rect -268 357 -246 359
rect -239 357 -234 359
rect -297 343 -256 345
rect -236 336 -234 357
rect -198 357 -196 389
rect -68 382 -66 395
rect -161 378 -159 380
rect -119 378 -117 381
rect -101 378 -99 381
rect -161 368 -159 372
rect -119 369 -117 373
rect -160 365 -159 368
rect -151 366 -117 369
rect -161 364 -159 365
rect -119 362 -117 366
rect -101 365 -99 373
rect -68 372 -66 376
rect -67 369 -66 372
rect -68 368 -66 369
rect -107 363 -99 365
rect -68 363 -66 365
rect -107 362 -106 363
rect -101 362 -99 363
rect -161 359 -159 361
rect -119 358 -117 359
rect -198 355 -166 357
rect -107 336 -106 359
rect -101 358 -99 359
rect -236 334 -106 336
rect -280 323 -231 325
rect -280 313 -278 323
rect -297 311 -274 313
rect -268 311 -267 313
rect -265 311 -246 313
rect -239 311 -236 313
rect -297 240 -295 311
rect -265 294 -263 311
rect -233 294 -231 323
rect -202 307 -200 309
rect -202 297 -200 301
rect -292 292 -274 294
rect -268 292 -263 294
rect -250 292 -246 294
rect -239 292 -231 294
rect -226 294 -206 297
rect -201 294 -200 297
rect -202 293 -200 294
rect -292 254 -290 292
rect -76 292 -74 305
rect -202 288 -200 290
rect -163 288 -161 290
rect -127 288 -125 291
rect -109 288 -107 291
rect -260 272 -256 275
rect -281 270 -274 272
rect -268 270 -246 272
rect -239 270 -234 272
rect -259 262 -257 270
rect -202 267 -200 284
rect -35 288 -33 291
rect -163 278 -161 282
rect -127 279 -125 283
rect -162 275 -161 278
rect -151 276 -125 279
rect -163 274 -161 275
rect -127 272 -125 276
rect -109 275 -107 283
rect -76 282 -74 286
rect -75 279 -74 282
rect -65 280 -52 283
rect -76 278 -74 279
rect -55 279 -52 280
rect -35 279 -33 283
rect -115 273 -107 275
rect -55 276 -33 279
rect -76 273 -74 275
rect -115 272 -114 273
rect -109 272 -107 273
rect -35 272 -33 276
rect -25 275 -23 304
rect 16 292 18 305
rect -17 288 -15 291
rect 63 287 65 289
rect 69 287 71 370
rect 73 287 75 289
rect 83 287 85 289
rect 93 287 95 289
rect 107 287 109 289
rect -17 275 -15 283
rect 16 282 18 286
rect 17 279 18 282
rect 16 278 18 279
rect 63 279 65 282
rect -25 273 -15 275
rect 69 279 71 282
rect 73 279 75 282
rect 83 280 85 282
rect 69 277 75 279
rect 16 273 18 275
rect -17 272 -15 273
rect 63 272 65 277
rect 73 272 75 277
rect 83 272 85 278
rect 93 280 95 282
rect 93 272 95 278
rect 107 277 109 282
rect 108 275 109 277
rect 107 272 109 275
rect -163 269 -161 271
rect -127 268 -125 269
rect -202 265 -168 267
rect -260 254 -256 259
rect -115 254 -114 269
rect -109 268 -107 269
rect -35 268 -33 269
rect -17 268 -15 269
rect 63 268 65 269
rect 73 268 75 269
rect 83 268 85 269
rect 93 268 95 269
rect 107 268 109 269
rect -292 252 -274 254
rect -268 252 -246 254
rect -239 252 -114 254
rect -297 238 -256 240
rect -280 210 -231 212
rect -280 200 -278 210
rect -297 198 -274 200
rect -268 198 -267 200
rect -265 198 -246 200
rect -239 198 -236 200
rect -297 127 -295 198
rect -265 181 -263 198
rect -233 181 -231 210
rect -109 202 -107 203
rect -95 202 -93 203
rect -79 202 -77 203
rect -65 202 -63 203
rect -50 202 -48 203
rect -21 202 -19 203
rect -202 194 -200 196
rect -165 194 -163 196
rect -109 190 -107 196
rect -202 184 -200 188
rect -165 184 -163 188
rect -108 187 -107 190
rect -95 188 -93 196
rect -79 188 -77 196
rect -65 188 -63 196
rect -50 188 -48 196
rect -21 192 -19 196
rect -292 179 -274 181
rect -268 179 -263 181
rect -250 179 -246 181
rect -239 179 -231 181
rect -226 181 -206 184
rect -201 181 -200 184
rect -164 181 -163 184
rect -109 182 -107 187
rect -95 182 -93 185
rect -79 182 -77 185
rect -65 182 -63 185
rect -50 182 -48 185
rect -21 182 -19 189
rect -202 180 -200 181
rect -165 180 -163 181
rect -292 141 -290 179
rect -202 175 -200 177
rect -109 178 -107 179
rect -95 178 -93 179
rect -79 178 -77 179
rect -65 178 -63 179
rect -50 178 -48 179
rect -21 178 -19 179
rect -165 175 -163 177
rect -196 171 -169 173
rect -165 171 -164 173
rect -260 159 -256 162
rect -281 157 -274 159
rect -268 157 -246 159
rect -239 157 -234 159
rect -254 150 -252 157
rect -260 145 -256 146
rect -260 142 -259 145
rect -257 142 -256 145
rect -260 141 -256 142
rect -292 139 -274 141
rect -268 139 -246 141
rect -239 139 -234 141
rect -297 125 -256 127
rect -280 66 -231 68
rect -280 56 -278 66
rect -297 54 -274 56
rect -268 54 -267 56
rect -265 54 -246 56
rect -239 54 -236 56
rect -297 -17 -295 54
rect -265 37 -263 54
rect -233 37 -231 66
rect -126 58 -124 59
rect -112 58 -110 59
rect -96 58 -94 59
rect -82 58 -80 59
rect -67 58 -65 59
rect -38 58 -36 59
rect -202 50 -200 52
rect -171 50 -169 52
rect -126 46 -124 52
rect -202 40 -200 44
rect -171 40 -169 44
rect -125 43 -124 46
rect -112 44 -110 52
rect -96 44 -94 52
rect -82 44 -80 52
rect -67 44 -65 52
rect -38 48 -36 52
rect -292 35 -274 37
rect -268 35 -263 37
rect -250 35 -246 37
rect -239 35 -231 37
rect -226 37 -206 40
rect -201 37 -200 40
rect -170 37 -169 40
rect -126 38 -124 43
rect -112 38 -110 41
rect -96 38 -94 41
rect -82 38 -80 41
rect -67 38 -65 41
rect -38 38 -36 45
rect -202 36 -200 37
rect -171 36 -169 37
rect -292 -3 -290 35
rect -202 31 -200 33
rect -126 34 -124 35
rect -112 34 -110 35
rect -96 34 -94 35
rect -82 34 -80 35
rect -67 34 -65 35
rect -38 34 -36 35
rect -171 31 -169 33
rect -260 15 -256 18
rect -281 13 -274 15
rect -268 13 -246 15
rect -239 13 -234 15
rect -254 7 -252 13
rect -260 1 -256 2
rect -260 -1 -259 1
rect -257 -1 -256 1
rect -260 -3 -256 -1
rect -292 -5 -274 -3
rect -268 -5 -246 -3
rect -239 -5 -234 -3
rect -297 -19 -256 -17
<< polycontact >>
rect -229 398 -226 402
rect -206 399 -201 402
rect -199 389 -196 391
rect -260 380 -256 384
rect -259 365 -257 367
rect -260 345 -256 349
rect -163 365 -160 368
rect -154 366 -151 369
rect -70 369 -67 372
rect 68 370 71 373
rect -166 355 -163 357
rect -229 293 -226 297
rect -206 294 -201 297
rect -25 304 -23 310
rect -202 284 -200 286
rect -260 275 -256 279
rect -165 275 -162 278
rect -156 276 -151 279
rect -78 279 -75 282
rect -69 280 -65 283
rect 14 279 17 282
rect 63 277 65 279
rect 82 278 85 280
rect 93 278 95 280
rect 107 275 108 277
rect -168 265 -163 267
rect -259 260 -257 262
rect -260 240 -256 244
rect -111 187 -108 190
rect -22 189 -19 192
rect -229 180 -226 184
rect -206 181 -201 184
rect -167 181 -164 184
rect -96 185 -93 188
rect -80 185 -77 188
rect -66 185 -63 188
rect -51 185 -48 188
rect -200 171 -196 173
rect -169 171 -165 173
rect -260 162 -256 166
rect -254 148 -252 150
rect -259 142 -257 145
rect -260 127 -256 131
rect -128 43 -125 46
rect -39 45 -36 48
rect -229 36 -226 40
rect -206 37 -201 40
rect -173 37 -170 40
rect -113 41 -110 44
rect -97 41 -94 44
rect -83 41 -80 44
rect -68 41 -65 44
rect -260 18 -256 22
rect -254 4 -252 7
rect -259 -1 -257 1
rect -260 -17 -256 -13
<< metal1 >>
rect -269 419 -245 423
rect -241 419 -221 423
rect -269 411 -245 415
rect -241 411 -226 415
rect -287 400 -273 404
rect -269 400 -245 404
rect -230 402 -226 411
rect -287 389 -283 400
rect -230 398 -229 402
rect -230 396 -226 398
rect -269 392 -245 396
rect -241 392 -226 396
rect -225 389 -221 419
rect -287 385 -262 389
rect -287 379 -273 383
rect -287 373 -283 375
rect -266 374 -262 385
rect -260 385 -221 389
rect -217 418 -185 420
rect -260 384 -256 385
rect -241 379 -228 383
rect -305 371 -283 373
rect -305 339 -303 371
rect -287 369 -283 371
rect -269 370 -245 374
rect -232 373 -228 375
rect -217 373 -214 418
rect -207 417 -203 418
rect -206 412 -203 417
rect -198 403 -195 408
rect -198 400 -191 403
rect -198 398 -195 400
rect -206 391 -203 394
rect -232 370 -214 373
rect -209 389 -199 391
rect -232 369 -228 370
rect -257 365 -254 367
rect -287 361 -273 365
rect -241 361 -228 365
rect -269 352 -245 356
rect -260 349 -256 352
rect -209 339 -207 389
rect -305 337 -207 339
rect -187 385 -185 418
rect -72 388 -61 389
rect -72 385 -69 388
rect -187 383 -69 385
rect -305 268 -303 337
rect -269 314 -245 318
rect -241 314 -221 318
rect -187 315 -185 383
rect -165 378 -162 383
rect -122 377 -120 383
rect -105 377 -103 383
rect -72 382 -69 383
rect -157 364 -154 374
rect -116 368 -114 374
rect -98 368 -96 375
rect -64 373 -61 378
rect -80 369 -70 372
rect -64 370 68 373
rect -80 368 -78 369
rect -116 366 -78 368
rect -64 368 -61 370
rect -98 362 -96 366
rect -165 357 -162 360
rect -72 361 -69 364
rect -122 357 -120 359
rect -72 359 -61 361
rect -72 357 -68 359
rect -163 355 -68 357
rect -269 306 -245 310
rect -241 306 -226 310
rect -287 295 -273 299
rect -269 295 -245 299
rect -230 297 -226 306
rect -287 284 -283 295
rect -230 293 -229 297
rect -230 291 -226 293
rect -269 287 -245 291
rect -241 287 -226 291
rect -225 284 -221 314
rect -287 280 -262 284
rect -287 274 -273 278
rect -287 268 -283 270
rect -266 269 -262 280
rect -260 280 -221 284
rect -217 313 -185 315
rect -260 279 -256 280
rect -241 274 -228 278
rect -305 266 -283 268
rect -305 234 -303 266
rect -287 264 -283 266
rect -269 265 -245 269
rect -232 268 -228 270
rect -217 268 -214 313
rect -207 312 -203 313
rect -206 307 -203 312
rect -198 298 -195 303
rect -198 295 -192 298
rect -187 295 -185 313
rect -25 310 -23 320
rect -80 298 -69 299
rect 12 298 61 300
rect -80 295 -77 298
rect 12 295 15 298
rect -198 293 -195 295
rect -187 293 15 295
rect -206 286 -203 289
rect -232 265 -214 268
rect -209 284 -202 286
rect -200 284 -196 286
rect -232 264 -228 265
rect -257 260 -254 262
rect -287 256 -273 260
rect -241 256 -228 260
rect -269 247 -245 251
rect -260 244 -256 247
rect -209 234 -207 284
rect -305 232 -207 234
rect -305 155 -303 232
rect -187 209 -185 293
rect -167 288 -164 293
rect -130 287 -128 293
rect -113 287 -111 293
rect -80 292 -77 293
rect -159 274 -156 284
rect -124 278 -122 284
rect -106 278 -104 285
rect -88 279 -78 282
rect -88 278 -86 279
rect -124 276 -86 278
rect -72 278 -69 288
rect -38 287 -36 293
rect -21 287 -19 293
rect 12 292 15 293
rect 59 292 61 298
rect -106 272 -104 276
rect -167 267 -164 270
rect -32 278 -30 284
rect -14 278 -12 285
rect 20 283 23 288
rect 59 290 109 292
rect 59 286 61 290
rect 104 286 106 290
rect 4 279 14 282
rect 20 280 43 283
rect 4 278 6 279
rect -32 276 6 278
rect 20 278 23 280
rect -80 271 -77 274
rect -14 272 -12 276
rect -130 267 -128 269
rect -80 269 -69 271
rect 41 279 43 280
rect 41 277 63 279
rect 96 277 98 283
rect 110 277 112 283
rect 66 275 107 277
rect 110 275 115 277
rect 12 271 15 274
rect 66 272 68 275
rect 76 272 78 275
rect 86 272 88 275
rect 96 272 98 275
rect 110 272 112 275
rect -80 267 -76 269
rect -38 267 -36 269
rect 12 269 23 271
rect 12 267 16 269
rect 59 267 61 270
rect 70 267 72 270
rect 80 267 82 270
rect 90 267 92 270
rect 104 267 106 270
rect -163 265 106 267
rect -187 206 -21 209
rect -269 201 -245 205
rect -241 201 -221 205
rect -187 202 -185 206
rect -269 193 -245 197
rect -241 193 -226 197
rect -287 182 -273 186
rect -269 182 -245 186
rect -230 184 -226 193
rect -287 171 -283 182
rect -230 180 -229 184
rect -230 178 -226 180
rect -269 174 -245 178
rect -241 174 -226 178
rect -225 171 -221 201
rect -287 167 -262 171
rect -287 161 -273 165
rect -287 155 -283 157
rect -266 156 -262 167
rect -260 167 -221 171
rect -217 201 -185 202
rect -113 201 -110 206
rect -217 200 -158 201
rect -260 166 -256 167
rect -241 161 -228 165
rect -305 153 -283 155
rect -305 121 -303 153
rect -287 151 -283 153
rect -269 152 -245 156
rect -232 155 -228 157
rect -217 155 -214 200
rect -207 199 -203 200
rect -206 194 -203 199
rect -187 199 -166 200
rect -198 180 -195 190
rect -206 173 -203 176
rect -232 152 -214 155
rect -209 171 -200 173
rect -232 151 -228 152
rect -287 143 -273 147
rect -254 146 -252 148
rect -241 143 -228 147
rect -269 134 -245 138
rect -260 131 -256 134
rect -209 121 -207 171
rect -305 119 -207 121
rect -305 11 -303 119
rect -187 65 -185 199
rect -169 194 -166 199
rect -99 201 -96 206
rect -83 201 -80 206
rect -106 192 -103 197
rect -69 201 -66 206
rect -92 192 -89 197
rect -55 201 -52 206
rect -76 192 -73 197
rect -25 202 -22 206
rect -62 192 -59 197
rect -47 192 -44 197
rect -18 192 -15 197
rect 79 192 81 231
rect -161 185 -158 190
rect -136 187 -111 190
rect -106 189 -22 192
rect -18 189 81 192
rect -136 185 -134 187
rect -69 185 -66 188
rect -161 182 -134 185
rect -44 182 -41 189
rect -18 182 -15 189
rect -161 180 -158 182
rect -169 173 -166 176
rect -113 174 -110 179
rect -25 174 -22 179
rect -113 173 -22 174
rect -170 171 -169 173
rect -165 171 -22 173
rect -187 62 -38 65
rect -269 57 -245 61
rect -241 57 -221 61
rect -187 58 -185 62
rect -269 49 -245 53
rect -241 49 -226 53
rect -287 38 -273 42
rect -269 38 -245 42
rect -230 40 -226 49
rect -287 27 -283 38
rect -230 36 -229 40
rect -230 34 -226 36
rect -269 30 -245 34
rect -241 30 -226 34
rect -225 27 -221 57
rect -287 23 -262 27
rect -287 17 -273 21
rect -287 11 -283 13
rect -266 12 -262 23
rect -260 23 -221 27
rect -217 56 -164 58
rect -130 57 -127 62
rect -260 22 -256 23
rect -241 17 -228 21
rect -305 9 -283 11
rect -305 -23 -303 9
rect -287 7 -283 9
rect -269 8 -245 12
rect -232 11 -228 13
rect -217 11 -214 56
rect -207 55 -203 56
rect -176 55 -172 56
rect -206 50 -203 55
rect -175 50 -172 55
rect -116 57 -113 62
rect -100 57 -97 62
rect -198 41 -195 46
rect -123 48 -120 53
rect -86 57 -83 62
rect -109 48 -106 53
rect -72 57 -69 62
rect -93 48 -90 53
rect -42 58 -39 62
rect -79 48 -76 53
rect -64 48 -61 53
rect -35 48 -32 53
rect 89 48 91 185
rect -167 41 -164 46
rect -146 43 -128 46
rect -123 45 -39 48
rect -35 45 91 48
rect -146 41 -144 43
rect -198 38 -192 41
rect -198 36 -195 38
rect -167 38 -144 41
rect -61 38 -58 45
rect -35 38 -32 45
rect -167 36 -164 38
rect -206 29 -203 32
rect -175 29 -172 32
rect -130 30 -127 35
rect -42 30 -39 35
rect -130 29 -39 30
rect -232 8 -214 11
rect -209 27 -39 29
rect -232 7 -228 8
rect -254 3 -252 4
rect -287 -1 -273 3
rect -241 -1 -228 3
rect -269 -10 -245 -6
rect -260 -13 -256 -10
rect -209 -23 -207 27
rect -305 -25 -207 -23
<< m2contact >>
rect -254 365 -252 367
rect -166 365 -163 368
rect -254 260 -251 262
rect -167 275 -165 278
rect 79 278 82 280
rect 91 278 93 280
rect 79 231 81 236
rect -254 142 -252 146
rect -259 140 -257 142
rect -99 185 -96 188
rect -169 181 -167 184
rect 89 185 91 191
rect -176 37 -173 40
rect -254 -2 -252 3
<< metal2 >>
rect -254 349 -252 365
rect -194 365 -166 368
rect -194 349 -192 365
rect -254 347 -192 349
rect -179 275 -167 278
rect -253 245 -251 260
rect -179 245 -177 275
rect -253 243 -177 245
rect 79 236 81 278
rect 89 191 91 280
rect -180 181 -169 184
rect -259 131 -257 140
rect -254 131 -252 142
rect -180 131 -178 181
rect -260 127 -256 131
rect -254 129 -178 131
rect -259 116 -257 127
rect -101 116 -99 188
rect -259 114 -99 116
rect -186 37 -176 40
rect -254 -13 -252 -2
rect -186 -13 -184 37
rect -254 -15 -184 -13
<< m123contact >>
rect -191 400 -189 403
rect -25 320 -23 325
rect -192 295 -189 298
rect -195 182 -192 185
rect -83 185 -80 188
rect -54 185 -51 188
rect -116 41 -113 44
rect -100 41 -97 44
rect -86 41 -83 44
rect -71 41 -68 44
rect -259 -4 -257 -1
<< metal3 >>
rect -191 327 -189 400
rect -191 325 -23 327
rect -191 238 -189 295
rect -191 236 -85 238
rect -87 188 -85 236
rect -51 219 -49 325
rect -59 217 -49 219
rect -59 188 -57 217
rect -87 185 -83 188
rect -59 185 -54 188
rect -192 182 -188 185
rect -190 79 -188 182
rect -87 79 -85 185
rect -190 77 -120 79
rect -122 44 -120 77
rect -106 77 -85 79
rect -106 44 -104 77
rect -59 74 -57 185
rect -89 72 -57 74
rect -89 44 -87 72
rect -122 41 -116 44
rect -106 41 -100 44
rect -89 41 -86 44
rect -76 41 -71 44
rect -259 -33 -257 -4
rect -76 -33 -74 41
rect -259 -35 -74 -33
<< labels >>
rlabel metal1 -246 -24 -246 -24 1 gnd
rlabel metal1 -215 56 -215 56 1 vdd
rlabel metal1 -193 40 -193 40 1 x0
rlabel polysilicon -258 15 -258 15 1 b0
rlabel polysilicon -258 -3 -258 -3 1 a0
rlabel polysilicon -258 142 -258 142 1 a1
rlabel polysilicon -259 159 -259 159 1 b1
rlabel m123contact -194 184 -194 184 1 x1
rlabel polysilicon -258 256 -258 256 1 a2
rlabel polysilicon -258 273 -258 273 1 b2
rlabel metal1 -193 297 -193 297 1 x2
rlabel polysilicon -258 360 -258 360 1 a3
rlabel polysilicon -258 379 -258 379 1 b3
rlabel metal1 -194 402 -194 402 1 x3
rlabel polycontact -155 278 -155 278 1 b2_not
rlabel metal1 -157 184 -157 184 1 b1_not
rlabel metal1 -164 39 -164 39 1 b0_not
rlabel metal1 -60 371 -60 371 1 AmoreB_3
rlabel metal1 24 281 24 281 1 AmoreB_2
rlabel metal1 -11 190 -11 190 1 AmoreB_1
rlabel metal1 -28 46 -28 46 1 AmoreB_0
rlabel metal1 113 276 113 276 7 out
rlabel metal1 -67 186 -67 186 1 temp
<< end >>
