* SPICE3 file created from final_4.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param width_P=8*LAMBDA
.param  width_N = 4*LAMBDA
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

* Vs0 s0 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
* Vs1 s1 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)

Vs0 s0 gnd DC 0
Vs1 s1 gnd DC 1.8

* Va3 a3 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
* Va2 a2 gnd PULSE(1.8 0 100ns 100ps 100ps 100ns 200ns)
* Va1 a1 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
* Va0 a0 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)

Va3 a3 gnd PULSE(0 1.8 0 100ps 100ps 200ns 400ns)
Va2 a2 gnd PULSE(0 1.8 0 100ps 100ps 200ns 400ns)
Va1 a1 gnd PULSE(0 1.8 0 100ps 100ps 200ns 400ns)
Va0 a0 gnd PULSE(0 1.8 0 100ps 100ps 200ns 400ns)

Vb3 b3 gnd DC 1.8
Vb2 b2 gnd DC 1.8
Vb1 b1 gnd DC 1.8
Vb0 b0 gnd DC 1.8

* Vb3 b3 gnd DC 1.8
* Vb2 b2 gnd DC 1.8
* Vb1 b1 gnd DC 1.8
* Vb0 b0 gnd DC 0

Vtempless temp_less gnd DC 1.8
Vtempmore temp_more gnd DC 1.8
Vtemp temp gnd DC 1.8
Vd2 equals_d gnd DC 1.8
* Vsmd smd gnd DC 1.8

.option scale=0.09u

M1000 adsub_b2 a_n33840_n2871# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=347733 ps=33048
M1001 a_n29457_n8883# a_n30123_n8919# vdd w_n29547_n8685# CMOSP w=54 l=18
+  ad=2916 pd=216 as=635202 ps=50436
M1002 a_n28620_n5877# x2 vdd w_n28737_n5787# CMOSP w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1003 gnd comp_a1 a_n30123_n1953# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1004 AlessB a_n27072_n891# vdd w_n27144_n792# CMOSP w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1005 gnd D1 a_n30483_5634# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1006 D1 a_n35820_n12033# gnd Gnd CMOSN w=27 l=18
+  ad=13122 pd=1026 as=0 ps=0
M1007 a_n29565_6714# a_n29286_7263# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1008 a_n33840_n1935# D gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1009 a_n28620_n1548# x2 vdd w_n28737_n1458# CMOSP w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1010 AmoreB_2 a_n27954_n5094# vdd w_n27576_n5085# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1011 comp_a0 comp_b0 a_n30123_n3051# w_n29898_n3420# CMOSP w=63 l=18
+  ad=6318 pd=450 as=6804 ps=468
M1012 comp_b0 a_n30330_n12609# a_n30123_n12177# Gnd CMOSN w=54 l=18
+  ad=7290 pd=594 as=5832 ps=432
M1013 D1 a_n30690_9612# a_n30483_10044# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=8748 ps=648
M1014 a_n29637_6840# a_n29853_7128# vdd w_n29718_6822# CMOSP w=45 l=18
+  ad=3240 pd=234 as=0 ps=0
M1015 AmoreB_3 a_n28710_n4284# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1016 a_n30123_n1953# a_n30330_n2187# a_n30123_n1755# w_n29898_n2124# CMOSP w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1017 a_n29673_7749# adsub_a2 a_n29673_7947# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=8748 ps=648
M1018 a_n30483_3897# adsub_a0 a_n29673_3897# w_n29448_3528# CMOSP w=63 l=18
+  ad=10206 pd=702 as=10206 ps=702
M1019 a_n33822_n15822# D3 vdd w_n33912_n15849# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1020 gnd comp_a3 a_n30330_n9351# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1021 a_n30123_n6282# comp_a1 a_n30123_n6084# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1022 comp_a2 a_n33822_n8721# vdd w_n33444_n8712# CMOSP w=54 l=18
+  ad=6318 pd=450 as=0 ps=0
M1023 a_n30483_7749# a_n30690_7515# a_n30483_7947# w_n30258_7578# CMOSP w=63 l=18
+  ad=6804 pd=468 as=10206 ps=702
M1024 a_n28773_n7326# b0_not gnd Gnd CMOSN w=27 l=18
+  ad=2916 pd=270 as=0 ps=0
M1025 a_n31851_n13896# and_a3 vdd w_n31941_n13923# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1026 a_n29286_5148# carry0 a_n29286_5022# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1027 a0_not comp_a0 vdd w_n29268_n2817# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1028 adsub_b3 a_n33840_n2376# vdd w_n33462_n2367# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1029 a_n33822_n8226# a3 vdd w_n33912_n8253# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1030 a_n31851_n14373# and_b2 vdd w_n31941_n14400# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1031 a_n33822_n14508# D3 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1032 adsub_a1 a_n33840_n1278# vdd w_n33462_n1269# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1033 a_n30123_n4320# comp_a3 a_n30123_n4122# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1034 a_n33822_n10638# D2 vdd w_n33912_n10665# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1035 and_b2 a_n33822_n14877# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1036 a_n33840_n2871# b2 vdd w_n33930_n2898# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1037 a_n30123_n5265# a_n30330_n5499# a_n30123_n5067# w_n29898_n5436# CMOSP w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1038 a_n35685_n12600# s1 a_n35820_n12600# Gnd CMOSN w=27 l=18
+  ad=243 pd=72 as=3159 ps=288
M1039 a_n28323_n5166# a_n28782_n5094# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1040 a_n28791_7749# carry1 sum2 Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1041 a_n33822_n8847# D2 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1042 a_n28224_n6030# temp_more a_n28350_n6030# Gnd CMOSN w=27 l=18
+  ad=3159 pd=288 as=2916 ps=270
M1043 a_n33822_n12573# D3 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1044 gnd D1 a_n30483_3699# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1045 a_n33822_n15291# b1 vdd w_n33912_n15318# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1046 a_n28782_n765# a2_not vdd w_n28872_n792# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1047 vdd adsub_a2 a_n29880_7515# w_n29448_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1048 gnd comp_a1 a_n30330_n6516# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1049 a_n29637_6723# a_n29853_7128# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1050 a_n30312_5085# adsub_a1 vdd w_n30402_5058# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1051 and_b1 a_n33822_n15291# vdd w_n33444_n15282# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1052 a3_not comp_a3 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1053 a_n30123_n7578# a_n30330_n7812# a_n30123_n7380# w_n29898_n7749# CMOSP w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1054 a_n27072_n5220# AmoreB_0 a_n26892_n5103# w_n27576_n5085# CMOSP w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1055 a_n29457_n9828# a_n30123_n9864# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1056 a_n28710_n4284# comp_a3 vdd w_n28800_n4311# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1057 a_n28152_n9981# a_n29457_n8883# gnd Gnd CMOSN w=27 l=18
+  ad=2916 pd=270 as=0 ps=0
M1058 a2_not comp_a2 vdd w_n29205_n675# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1059 x1 a_n30123_n6084# vdd w_n29547_n5850# CMOSP w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1060 a_n30123_n12375# comp_a0 a_n30123_n12177# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1061 a_n33822_n9135# D2 vdd w_n33912_n9162# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1062 a_n34407_n1233# D1 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1063 a_n35820_n12888# s0 a_n35703_n13014# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=729 ps=108
M1064 comp_b2 comp_a2 a_n30123_n9864# w_n29898_n10233# CMOSP w=63 l=18
+  ad=9720 pd=684 as=6804 ps=468
M1065 vdd comp_a2 a_n30330_n5499# w_n29898_n5436# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1066 D0 a_n35820_n11565# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1067 x1 a_n30123_n1755# vdd w_n29547_n1521# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1068 a_n35820_n12033# s1_not a_n35820_n12159# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1069 x3 a_n30123_n4122# vdd w_n29547_n3888# CMOSP w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1070 vdd comp_b2 a_n30330_n1170# w_n29898_n1107# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1071 a_n27756_n9981# a_n29457_n12141# a_n27882_n9981# Gnd CMOSN w=27 l=18
+  ad=3159 pd=288 as=2916 ps=270
M1072 a_n26892_n774# AlessB_1 a_n26982_n774# w_n27144_n792# CMOSP w=45 l=18
+  ad=3240 pd=234 as=3240 ps=234
M1073 a_n28791_9846# a_n28998_9612# sum3 w_n28566_9675# CMOSP w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1074 vdd a_n30285_n7686# a_n30330_n7812# w_n29898_n7749# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1075 comp_b0 comp_a0 a_n30123_n12177# w_n29898_n12546# CMOSP w=63 l=18
+  ad=9720 pd=684 as=6804 ps=468
M1076 comp_a0 a_n33822_n9666# gnd Gnd CMOSN w=27 l=18
+  ad=4374 pd=378 as=0 ps=0
M1077 vdd carry0 a_n28998_5400# w_n28566_5463# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1078 a_n30483_9846# a_n30690_9612# a_n30483_10044# w_n30258_9675# CMOSP w=63 l=18
+  ad=6804 pd=468 as=10206 ps=702
M1079 a_n33840_n864# D vdd w_n33930_n891# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1080 a_n33822_n11709# D2 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1081 a_n26811_n9945# k gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1082 vdd comp_b0 a_n30330_n3483# w_n29898_n3420# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1083 gnd comp_a0 a_n30330_n12609# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1084 a_n33822_n13887# a0 a_n33822_n14013# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1085 a_n28683_n891# comp_b2 a_n28782_n891# Gnd CMOSN w=27 l=9
+  ad=1215 pd=144 as=2430 ps=234
M1086 vdd D1 a_n28998_3465# w_n28566_3528# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1087 a_n33840_n3816# b0 a_n33840_n3942# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1088 a_n33822_n10143# b3 vdd w_n33912_n10170# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1089 gnd comp_a3 a_n30330_n4554# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1090 a_n30312_3150# adsub_a0 vdd w_n30402_3123# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1091 a_n28503_n2997# x2 a_n28647_n2997# Gnd CMOSN w=27 l=18
+  ad=2916 pd=270 as=3402 ps=306
M1092 comp_b3 a_n33822_n10143# vdd w_n33444_n10134# CMOSP w=54 l=18
+  ad=9720 pd=684 as=0 ps=0
M1093 a_n26892_n5103# AmoreB_1 a_n26982_n5103# w_n27576_n5085# CMOSP w=45 l=18
+  ad=0 pd=0 as=3240 ps=234
M1094 a_n31851_n13896# and_b3 vdd w_n31941_n13923# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1095 a_n30123_n9117# a_n30330_n9351# a_n30123_n8919# w_n29898_n9288# CMOSP w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1096 vdd a_n29673_10044# a_n28791_9846# w_n28566_9675# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1097 gnd adsub_a1 a_n29880_5400# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1098 a_n31851_n15237# and_a0 vdd w_n31941_n15264# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1099 a_n28377_n7326# x3 a_n28503_n7326# Gnd CMOSN w=27 l=18
+  ad=3159 pd=288 as=2916 ps=270
M1100 b0_not comp_b0 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1101 b1_not comp_b1 vdd w_n29214_n5850# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1102 a_n27072_n5220# AmoreB_3 gnd Gnd CMOSN w=27 l=18
+  ad=2916 pd=432 as=0 ps=0
M1103 a_n29637_8820# a_n29565_8811# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1104 a_n34407_n1233# D0 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1105 a_n33822_n12447# a3 vdd w_n33912_n12474# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1106 a_n28152_n9828# a_n29457_n9828# vdd w_n28260_n9846# CMOSP w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1107 a_n28773_n7173# b0_not vdd w_n28890_n7083# CMOSP w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1108 a_n28791_5634# a_n28998_5400# sum1 w_n28566_5463# CMOSP w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1109 and_oper_out2 a_n31851_n14373# vdd w_n31473_n14364# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1110 a0_not comp_a0 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1111 a_n33822_n14382# D3 vdd w_n33912_n14409# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1112 a1_not comp_a1 vdd w_n29214_n1521# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1113 gnd adsub_a0 a_n29880_3465# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1114 a_n30123_9# comp_b3 a_n30123_207# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1115 a_n33840_n369# a3 a_n33840_n495# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1116 a_n33840_n1809# a0 a_n33840_n1935# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1117 a_n33840_n2502# D gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1118 and_a3 a_n33822_n12447# vdd w_n33444_n12438# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1119 vdd adsub_b1 a_n30690_5400# w_n30258_5463# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1120 a_n33822_n11052# b1 a_n33822_n11178# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1121 gnd a_n30483_10044# a_n29673_9846# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1122 a_n27954_n765# x3 vdd w_n28044_n792# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1123 a_n29853_3078# a_n30312_3150# vdd w_n29934_3159# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1124 a_n30483_7947# adsub_a2 a_n29673_7947# w_n29448_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=10206 ps=702
M1125 vdd adsub_b0 a_n30690_3465# w_n30258_3528# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1126 a_n33822_n13068# D3 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1127 a_n29673_5634# adsub_a1 a_n29673_5832# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=8748 ps=648
M1128 a_n30312_3150# adsub_a0 a_n30312_3024# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1129 gnd carry0 a_n28998_5400# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1130 a_n28620_n5877# b1_not vdd w_n28737_n5787# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1131 vdd D1 a_n30483_9846# w_n30258_9675# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1132 a_n27954_n5094# x3 a_n27954_n5220# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1133 a_n30123_n12375# a_n30330_n12609# a_n30123_n12177# w_n29898_n12546# CMOSP w=63 l=18
+  ad=6804 pd=468 as=0 ps=0
M1134 a_n31851_n14022# and_a3 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1135 a_n28620_n1548# a1_not vdd w_n28737_n1458# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1136 b2_not comp_b2 vdd w_n29205_n5004# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1137 a_n28782_n765# comp_b2 vdd w_n28872_n792# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1138 a_n30483_5634# a_n30690_5400# a_n30483_5832# w_n30258_5463# CMOSP w=63 l=18
+  ad=6804 pd=468 as=10206 ps=702
M1139 x1 a_n30123_n6084# gnd Gnd CMOSN w=27 l=18
+  ad=2916 pd=324 as=0 ps=0
M1140 gnd D1 a_n28998_3465# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1141 gnd adsub_b3 a_n30690_9612# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1142 comp_b2 a_n30330_n5499# a_n30123_n5067# Gnd CMOSN w=54 l=18
+  ad=7290 pd=594 as=5832 ps=432
M1143 gnd a_n29673_10044# a_n28791_9846# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1144 a_n29286_5148# carry0 vdd w_n29376_5121# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1145 vdd comp_b3 a_n30123_n9117# w_n29898_n9288# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1146 adsub_a0 a_n33840_n1809# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1147 k a_n28152_n9828# gnd Gnd CMOSN w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
M1148 a_n33822_n8721# a2 a_n33822_n8847# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1149 a_n28791_3699# a_n28998_3465# sum0 w_n28566_3528# CMOSP w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1150 a_n28620_n5877# x3 a_n28224_n6030# Gnd CMOSN w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1151 a_n29286_5022# a_n29673_5832# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1152 a_n29853_3078# a_n30312_3150# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1153 a_n35820_n12888# s1 vdd w_n35910_n12915# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1154 a_n33822_n8721# D2 vdd w_n33912_n8748# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1155 x3 a_n30123_n4122# gnd Gnd CMOSN w=27 l=18
+  ad=2916 pd=324 as=0 ps=0
M1156 a_n28791_5634# carry0 sum1 Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1157 a_n29673_5832# carry0 sum1 w_n28566_5463# CMOSP w=63 l=18
+  ad=10206 pd=702 as=0 ps=0
M1158 vdd comp_a0 a_n30330_n12609# w_n29898_n12546# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1159 carry1 a_n29637_4608# vdd w_n29718_4707# CMOSP w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1160 a_n27018_n5103# AmoreB_3 a_n27072_n5103# w_n27576_n5085# CMOSP w=45 l=18
+  ad=810 pd=126 as=1620 ps=162
M1161 and_oper_out1 a_n31851_n14769# vdd w_n31473_n14760# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1162 comp_a0 a_n30330_n3483# a_n30123_n3051# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1163 a_n33822_n11583# D2 vdd w_n33912_n11610# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1164 adsub_b1 a_n33840_n3285# vdd w_n33462_n3276# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1165 and_b0 a_n33822_n15822# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1166 a_n33822_n9135# a1 vdd w_n33912_n9162# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1167 a_n30483_10044# a_n29880_9612# a_n29673_10044# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=8748 ps=648
M1168 a_n31851_n14769# and_a1 vdd w_n31941_n14796# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1169 a_n33822_n15417# D3 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1170 a_n30123_n11079# comp_a1 a_n30123_n10881# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1171 a_n29673_3699# adsub_a0 a_n29673_3897# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=8748 ps=648
M1172 a_n30123_n1953# comp_b1 a_n30123_n1755# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1173 a_n30312_5085# a_n30483_5832# vdd w_n30402_5058# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1174 carry0 a_n29637_2673# vdd w_n29718_2772# CMOSP w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1175 a_n31851_n15237# and_b0 vdd w_n31941_n15264# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1176 a_n33822_n9792# D2 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1177 a_n28494_n6030# comp_a1 a_n28620_n6030# Gnd CMOSN w=27 l=18
+  ad=3402 pd=306 as=2916 ps=270
M1178 comp_a3 a_n33822_n8226# gnd Gnd CMOSN w=27 l=18
+  ad=4374 pd=378 as=0 ps=0
M1179 AlessB_0 a_n28773_n2844# gnd Gnd CMOSN w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
M1180 and_oper_out3 a_n31851_n13896# vdd w_n31473_n13887# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1181 gnd comp_b3 a_n30330_n225# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1182 a_n33822_n13482# D3 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1183 a_n30483_5832# a_n29880_5400# a_n29673_5832# Gnd CMOSN w=54 l=18
+  ad=8748 pd=648 as=0 ps=0
M1184 a_n33822_n13887# D3 vdd w_n33912_n13914# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1185 a_n33822_n10269# D2 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1186 a_n30483_3699# a_n30690_3465# a_n30483_3897# w_n30258_3528# CMOSP w=63 l=18
+  ad=6804 pd=468 as=0 ps=0
M1187 a_n28152_n9828# temp a_n27756_n9981# Gnd CMOSN w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1188 a_n28773_n7173# x3 vdd w_n28890_n7083# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1189 a_n35820_n12033# s1_not vdd w_n35910_n12060# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1190 b1_not comp_b1 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1191 gnd D1 a_n30483_7749# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1192 a_n35820_n11691# s0_not gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1193 D1 adsub_b1 a_n30483_5832# w_n30258_5463# CMOSP w=63 l=18
+  ad=16524 pd=1152 as=0 ps=0
M1194 a_n29286_3213# D1 vdd w_n29376_3186# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1195 a_n28224_n1701# temp_less a_n28350_n1701# Gnd CMOSN w=27 l=18
+  ad=3159 pd=288 as=2916 ps=270
M1196 a_n29286_3213# D1 a_n29286_3087# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1197 a_n26811_n9819# equals_d a_n26811_n9945# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1198 carry1 a_n29637_4608# gnd Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1199 a_n30123_n5265# comp_a2 a_n30123_n5067# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1200 a_n28791_3699# D1 sum0 Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1201 a_n29637_8820# a_n29853_9225# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1202 a_n29673_3897# D1 sum0 w_n28566_3528# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1203 D2 a_n35820_n12474# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1204 AlessB_2 a_n27954_n765# vdd w_n27576_n756# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1205 adsub_a3 a_n33840_n369# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1206 carry0 a_n29637_2673# gnd Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1207 adsub_a2 a_n33840_n864# vdd w_n33462_n855# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1208 a_n29673_5832# a_n28998_5400# sum1 Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1209 vdd comp_b1 a_n30123_n6282# w_n29898_n6453# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1210 a_n31851_n13896# and_b3 a_n31851_n14022# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1211 a_n30123_n7578# a_n30285_n7686# a_n30123_n7380# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1212 a_n33822_n10638# b2 a_n33822_n10764# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1213 a_n28773_n2844# x2 vdd w_n28890_n2754# CMOSP w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1214 a_n28773_n7173# a_n30285_n7686# a_n28377_n7326# Gnd CMOSN w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1215 a_n27954_n5094# x3 vdd w_n28044_n5121# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1216 vdd a_n30483_5832# a_n29673_5634# w_n29448_5463# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1217 a_n26982_n5103# AmoreB_3 a_n27018_n5103# w_n27576_n5085# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1218 a_n30312_3150# a_n30483_3897# vdd w_n30402_3123# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1219 gnd comp_b1 a_n30123_n11079# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1220 a_n29673_10044# a_n28998_9612# sum3 Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1221 comp_a2 a_n30330_n1170# a_n30123_n738# Gnd CMOSN w=54 l=18
+  ad=4374 pd=378 as=5832 ps=432
M1222 a_n33840_n2376# b3 a_n33840_n2502# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1223 comp_b2 a_n33822_n10638# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1224 a_n28323_n837# a_n28782_n765# vdd w_n28404_n756# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1225 a_n30483_3897# a_n29880_3465# a_n29673_3897# Gnd CMOSN w=54 l=18
+  ad=8748 pd=648 as=0 ps=0
M1226 a_n29457_n12141# a_n30123_n12177# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1227 comp_b2 a_n30330_n10296# a_n30123_n9864# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1228 AmoreB_1 a_n28620_n5877# vdd w_n28737_n5787# CMOSP w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1229 gnd comp_a2 a_n30330_n5499# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1230 vdd comp_b3 a_n30123_n4320# w_n29898_n4491# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1231 a_n29637_8820# a_n29565_8811# a_n29637_8937# w_n29718_8919# CMOSP w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1232 a_n33822_n11052# b1 vdd w_n33912_n11079# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1233 gnd comp_a2 a_n30330_n10296# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1234 AlessB_1 a_n28620_n1548# vdd w_n28737_n1458# CMOSP w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1235 gnd comp_b2 a_n30330_n1170# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1236 comp_a2 comp_b2 a_n30123_n738# w_n29898_n1107# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1237 AequalsB a_n26811_n9819# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1238 a_n28647_n7326# x1 a_n28773_n7326# Gnd CMOSN w=27 l=18
+  ad=3402 pd=306 as=0 ps=0
M1239 comp_b1 a_n33822_n11052# vdd w_n33444_n11043# CMOSP w=54 l=18
+  ad=9720 pd=684 as=0 ps=0
M1240 a_n30483_7749# adsub_b2 a_n30483_7947# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=8748 ps=648
M1241 vdd carry1 a_n28998_7515# w_n28566_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1242 a_n30312_7200# adsub_a2 vdd w_n30402_7173# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1243 a_n33840_n495# D gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1244 D1 adsub_b0 a_n30483_3897# w_n30258_3528# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1245 a_n30312_7200# adsub_a2 a_n30312_7074# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1246 gnd a_n30285_n7686# a_n30330_n7812# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1247 x2 a_n30123_n5067# vdd w_n29547_n4833# CMOSP w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1248 a_n30123_9# a_n30330_n225# a_n30123_207# w_n29898_n162# CMOSP w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1249 AlessB_3 a_n28710_45# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1250 a_n31851_n14769# and_b1 vdd w_n31941_n14796# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1251 a_n30123_n11079# a_n30330_n11313# a_n30123_n10881# w_n29898_n11250# CMOSP w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1252 a_n27954_n891# a_n28323_n837# gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1253 a_n33822_n13356# a1 vdd w_n33912_n13383# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1254 a_n29673_9846# a_n29880_9612# a_n29673_10044# w_n29448_9675# CMOSP w=63 l=18
+  ad=6804 pd=468 as=10206 ps=702
M1255 gnd comp_a2 a_n30123_n936# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1256 gnd comp_b0 a_n30330_n3483# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1257 a_n27018_n774# AlessB_3 a_n27072_n774# w_n27144_n792# CMOSP w=45 l=18
+  ad=810 pd=126 as=1620 ps=162
M1258 a_n33822_n15291# D3 vdd w_n33912_n15318# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1259 a_n33840_n3411# D gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1260 and_a1 a_n33822_n13356# vdd w_n33444_n13347# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1261 a_n33840_n3816# D vdd w_n33930_n3843# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1262 a_n30312_3024# a_n30483_3897# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1263 a_n35820_n11565# s1_not vdd w_n35910_n11592# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1264 a_n29673_3897# a_n28998_3465# sum0 Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1265 x2 a_n30123_n738# gnd Gnd CMOSN w=27 l=18
+  ad=2916 pd=324 as=0 ps=0
M1266 and_oper_out0 a_n31851_n15237# vdd w_n31473_n15228# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1267 gnd adsub_a2 a_n29880_7515# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1268 vdd a_n30483_3897# a_n29673_3699# w_n29448_3528# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1269 AlessB_3 a_n28710_45# vdd w_n28332_54# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1270 a_n28710_45# comp_b3 a_n28611_n81# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=1215 ps=144
M1271 vdd comp_a2 a_n30123_n936# w_n29898_n1107# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1272 a_n30123_n9117# comp_a3 a_n30123_n8919# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1273 adsub_b2 a_n33840_n2871# vdd w_n33462_n2862# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1274 a_n28350_n6030# x2 a_n28494_n6030# Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1275 x0 a_n30123_n3051# vdd w_n29547_n2817# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1276 a_n33822_n8721# a2 vdd w_n33912_n8748# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1277 a_n29853_7128# a_n30312_7200# vdd w_n29934_7209# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1278 D1 a_n35820_n12033# vdd w_n35442_n12024# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1279 a_n35820_n13014# s1 gnd Gnd CMOSN w=27 l=18
+  ad=2673 pd=252 as=0 ps=0
M1280 vdd adsub_b2 a_n30690_7515# w_n30258_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1281 a_n33840_n1404# D gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1282 D a_n34407_n1233# gnd Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1283 a_n33840_n1809# D vdd w_n33930_n1836# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1284 a_n29286_5148# a_n29673_5832# vdd w_n29376_5121# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1285 a_n28611_n4410# comp_a3 a_n28710_n4410# Gnd CMOSN w=27 l=9
+  ad=1215 pd=144 as=2430 ps=234
M1286 a_n35820_n12159# s0 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1287 AmoreB_3 a_n28710_n4284# vdd w_n28332_n4275# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1288 a_n35820_n12474# s1 a_n35685_n12600# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1289 a_n29565_8811# a_n29286_9360# vdd w_n28908_9369# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1290 a_n33822_n9666# a0 a_n33822_n9792# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1291 gnd carry1 a_n28998_7515# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1292 adsub_b0 a_n33840_n3816# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1293 s0_not s0 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1294 vdd comp_b1 a_n30123_n11079# w_n29898_n11250# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1295 a_n27882_n9981# a_n29457_n10845# a_n28026_n9981# Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=3402 ps=306
M1296 a_n33822_n14013# D3 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1297 a_n33822_n14877# b2 vdd w_n33912_n14904# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1298 AlessB_0 a_n28773_n2844# vdd w_n28890_n2754# CMOSP w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1299 a_n28773_n7173# a_n30285_n7686# vdd w_n28890_n7083# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1300 a_n33822_n10143# D2 vdd w_n33912_n10170# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1301 a_n29853_7128# a_n30312_7200# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1302 and_b3 a_n33822_n14382# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1303 a3_not comp_a3 vdd w_n29178_135# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1304 and_b2 a_n33822_n14877# vdd w_n33444_n14868# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1305 a_n30483_9846# adsub_b3 a_n30483_10044# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1306 a_n28773_n2997# a0_not gnd Gnd CMOSN w=27 l=18
+  ad=2916 pd=270 as=0 ps=0
M1307 a_n29286_7263# carry1 vdd w_n29376_7236# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1308 vdd comp_a2 a_n30330_n10296# w_n29898_n10233# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1309 a_n33822_n8352# D2 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1310 a_n28323_n5166# a_n28782_n5094# vdd w_n28404_n5085# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1311 a_n28620_n1548# x3 a_n28224_n1701# Gnd CMOSN w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1312 s1_not s1 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1313 vdd comp_b3 a_n30330_n225# w_n29898_n162# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1314 gnd comp_b3 a_n30123_n9117# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1315 a_n33822_n12447# D3 vdd w_n33912_n12474# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1316 a_n29565_8811# a_n29286_9360# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1317 a_n29673_7947# carry1 sum2 w_n28566_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1318 carry2 a_n29637_6723# vdd w_n29718_6822# CMOSP w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1319 a_n29286_3213# a_n29673_3897# vdd w_n29376_3186# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1320 a_n28773_n7173# x1 vdd w_n28890_n7083# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1321 a_n27954_n5220# a_n28323_n5166# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1322 a_n29457_n9828# a_n30123_n9864# vdd w_n29547_n9630# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1323 a_n29286_3087# a_n29673_3897# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1324 a_n33822_n11178# D2 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1325 x2 a_n30123_n5067# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1326 a_n29637_8937# a_n29853_9225# vdd w_n29718_8919# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1327 gnd adsub_b1 a_n30690_5400# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1328 a_n28152_n9828# a_n29457_n8883# vdd w_n28260_n9846# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1329 a_n34407_n1233# D1 a_n34407_n1116# w_n34488_n1134# CMOSP w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1330 comp_b2 a_n33822_n10638# vdd w_n33444_n10629# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1331 a_n30123_n3249# a_n30330_n3483# a_n30123_n3051# w_n29898_n3420# CMOSP w=63 l=18
+  ad=6804 pd=468 as=0 ps=0
M1332 a_n28494_n1701# comp_b1 a_n28620_n1701# Gnd CMOSN w=27 l=18
+  ad=3402 pd=306 as=2916 ps=270
M1333 D0 a_n35820_n11565# vdd w_n35442_n11556# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1334 a_n29457_n10845# a_n30123_n10881# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1335 b3_not comp_b3 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1336 a_n29457_n7344# a_n30123_n7380# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1337 gnd adsub_b0 a_n30690_3465# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1338 a_n27072_n891# AlessB_3 gnd Gnd CMOSN w=27 l=18
+  ad=2916 pd=432 as=0 ps=0
M1339 a_n30483_7947# a_n29880_7515# a_n29673_7947# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1340 a_n33822_n12942# a2 vdd w_n33912_n12969# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1341 a_n29286_7263# carry1 a_n29286_7137# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1342 x0 a_n30123_n3051# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1343 and_a2 a_n33822_n12942# vdd w_n33444_n12933# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1344 gnd D1 a_n30483_9846# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1345 a_n28152_n9828# a_n29457_n12141# vdd w_n28260_n9846# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1346 comp_b0 a_n30285_n7686# a_n30123_n7380# w_n29898_n7749# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1347 comp_a0 a_n33822_n9666# vdd w_n33444_n9657# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1348 a_n33822_n15822# b0 a_n33822_n15948# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1349 comp_a1 a_n33822_n9135# gnd Gnd CMOSN w=27 l=18
+  ad=4374 pd=378 as=0 ps=0
M1350 D1 adsub_b2 a_n30483_7947# w_n30258_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1351 a_n33840_n2376# D vdd w_n33930_n2403# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1352 carry2 a_n29637_6723# gnd Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1353 a_n30483_5634# adsub_b1 a_n30483_5832# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1354 comp_b0 a_n33822_n11583# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1355 a_n26811_n9819# k vdd w_n26901_n9846# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1356 vdd adsub_a3 a_n29880_9612# w_n29448_9675# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1357 a_n33840_n3285# b1 a_n33840_n3411# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1358 a_n27072_n891# AlessB_0 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1359 a_n33840_n3816# b0 vdd w_n33930_n3843# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1360 a_n30312_7200# a_n30483_7947# vdd w_n30402_7173# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1361 a_n27072_n891# AlessB_2 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1362 a_n30312_7074# a_n30483_7947# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1363 a_n29673_7947# a_n28998_7515# sum2 Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1364 b0_not comp_b0 vdd w_n29268_n7146# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1365 and_a0 a_n33822_n13887# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1366 gnd comp_b1 a_n30123_n6282# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1367 a_n34407_n1116# D0 vdd w_n34488_n1134# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1368 a_n28683_n5220# comp_a2 a_n28782_n5220# Gnd CMOSN w=27 l=9
+  ad=1215 pd=144 as=2430 ps=234
M1369 a_n33840_n1278# a1 a_n33840_n1404# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1370 a_n28377_n2997# x3 a_n28503_n2997# Gnd CMOSN w=27 l=18
+  ad=3159 pd=288 as=0 ps=0
M1371 a_n33840_n369# a3 vdd w_n33930_n396# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1372 a_n33840_n1809# a0 vdd w_n33930_n1836# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1373 vdd comp_a0 a_n30123_n3249# w_n29898_n3420# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1374 AlessB a_n27072_n891# gnd Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1375 a_n29457_n8883# a_n30123_n8919# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1376 gnd comp_b3 a_n30123_n4320# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1377 x3 a_n30123_207# vdd w_n29547_441# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1378 vdd comp_b1 a_n30330_n2187# w_n29898_n2124# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1379 a_n30312_5085# adsub_a1 a_n30312_4959# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1380 a_n28710_n81# a3_not gnd Gnd CMOSN w=27 l=18
+  ad=2430 pd=234 as=0 ps=0
M1381 a_n35820_n12033# s0 vdd w_n35910_n12060# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1382 a_n35820_n12474# s1 vdd w_n35910_n12501# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1383 AmoreB_2 a_n27954_n5094# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1384 vdd comp_b2 a_n30123_n5265# w_n29898_n5436# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1385 comp_b3 comp_a3 a_n30123_n8919# w_n29898_n9288# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1386 a_n28620_n6030# b1_not gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1387 a_n30483_3699# adsub_b0 a_n30483_3897# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1388 a_n30312_9297# adsub_a3 a_n30312_9171# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1389 a_n28782_n5220# b2_not gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1390 a_n27954_n5094# a_n28323_n5166# vdd w_n28044_n5121# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1391 vdd a_n30483_7947# a_n29673_7749# w_n29448_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1392 vdd comp_b0 a_n30123_n7578# w_n29898_n7749# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1393 D1 a_n30690_5400# a_n30483_5832# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1394 vdd a_n29673_5832# a_n28791_5634# w_n28566_5463# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1395 a_n33822_n14877# b2 a_n33822_n15003# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1396 a_n29637_4608# a_n29565_4599# a_n29637_4725# w_n29718_4707# CMOSP w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1397 comp_a2 a_n33822_n8721# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1398 a_n28611_n81# comp_b3 a_n28710_n81# Gnd CMOSN w=27 l=9
+  ad=0 pd=0 as=0 ps=0
M1399 a_n33822_n8226# a3 a_n33822_n8352# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1400 gnd comp_b0 a_n30123_n12375# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1401 adsub_b3 a_n33840_n2376# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1402 D3 a_n35820_n12888# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1403 a_n28350_n1701# x2 a_n28494_n1701# Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1404 adsub_a0 a_n33840_n1809# vdd w_n33462_n1800# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1405 a_n33822_n10764# D2 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1406 x3 a_n30123_207# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1407 a_n28773_n2844# a0_not vdd w_n28890_n2754# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1408 a_n29637_2673# a_n29565_2664# a_n29637_2790# w_n29718_2772# CMOSP w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1409 a_n29853_9225# a_n30312_9297# vdd w_n29934_9306# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1410 k a_n28152_n9828# vdd w_n28260_n9846# CMOSP w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1411 a_n30123_n10062# a_n30330_n10296# a_n30123_n9864# w_n29898_n10233# CMOSP w=63 l=18
+  ad=6804 pd=468 as=0 ps=0
M1412 a_n28782_n891# a2_not gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1413 gnd a_n30483_5832# a_n29673_5634# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1414 and_a2 a_n33822_n12942# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1415 a_n27072_n5220# AmoreB_2 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1416 a_n28620_n5877# temp_more vdd w_n28737_n5787# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1417 a_n29286_7263# a_n29673_7947# vdd w_n29376_7236# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1418 a_n29673_10044# carry2 sum3 w_n28566_9675# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1419 a_n28782_n5094# comp_a2 a_n28683_n5220# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1420 and_b0 a_n33822_n15822# vdd w_n33444_n15813# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1421 a_n33822_n11052# D2 vdd w_n33912_n11079# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1422 and_b1 a_n33822_n15291# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1423 a_n28620_n1548# temp_less vdd w_n28737_n1458# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1424 vdd D1 a_n30483_5634# w_n30258_5463# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1425 a2_not comp_a2 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1426 D1 adsub_b3 a_n30483_10044# w_n30258_9675# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1427 vdd comp_a3 a_n30123_9# w_n29898_n162# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1428 comp_a3 a_n33822_n8226# vdd w_n33444_n8217# CMOSP w=54 l=18
+  ad=6318 pd=450 as=0 ps=0
M1429 a_n33822_n9261# D2 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1430 a_n29637_4608# a_n29565_4599# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1431 a_n33822_n9666# D2 vdd w_n33912_n9693# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1432 AmoreB a_n27072_n5220# gnd Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1433 D1 a_n30690_3465# a_n30483_3897# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1434 a_n33822_n13356# D3 vdd w_n33912_n13383# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1435 vdd a_n29673_3897# a_n28791_3699# w_n28566_3528# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1436 a_n29673_7749# a_n29880_7515# a_n29673_7947# w_n29448_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1437 x1 a_n30123_n1755# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1438 gnd a_n29673_5832# a_n28791_5634# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1439 a_n29637_2673# a_n29565_2664# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1440 comp_b1 comp_a1 a_n30123_n6084# w_n29898_n6453# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1441 a_n29853_9225# a_n30312_9297# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1442 a_n33840_n2376# b3 vdd w_n33930_n2403# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1443 a_n28152_n9828# temp vdd w_n28260_n9846# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1444 a_n35820_n11565# s0_not vdd w_n35910_n11592# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1445 a_n27072_n891# AlessB_1 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1446 a_n33822_n15822# b0 vdd w_n33912_n15849# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1447 a_n29286_9360# carry2 vdd w_n29376_9333# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1448 a_n29565_4599# a_n29286_5148# vdd w_n28908_5157# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1449 comp_b1 a_n30330_n11313# a_n30123_n10881# Gnd CMOSN w=54 l=18
+  ad=7290 pd=594 as=0 ps=0
M1450 comp_a1 comp_b1 a_n30123_n1755# w_n29898_n2124# CMOSP w=63 l=18
+  ad=6318 pd=450 as=0 ps=0
M1451 a_n29673_9846# adsub_a3 a_n29673_10044# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1452 a_n29286_7137# a_n29673_7947# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1453 a_n26811_n9819# equals_d vdd w_n26901_n9846# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1454 a_n33840_n2997# D gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1455 a_n28503_n7326# x2 a_n28647_n7326# Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1456 gnd a_n30483_3897# a_n29673_3699# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1457 comp_a3 a_n30330_n225# a_n30123_207# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1458 comp_b3 comp_a3 a_n30123_n4122# w_n29898_n4491# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1459 D2 a_n35820_n12474# vdd w_n35442_n12465# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1460 adsub_a3 a_n33840_n369# vdd w_n33462_n360# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1461 a_n33822_n14382# b3 a_n33822_n14508# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1462 a_n28782_n5094# b2_not vdd w_n28872_n5121# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1463 gnd adsub_b2 a_n30690_7515# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1464 a_n33822_n10638# b2 vdd w_n33912_n10665# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1465 vdd D1 a_n30483_3699# w_n30258_3528# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1466 comp_b3 a_n33822_n10143# gnd Gnd CMOSN w=27 l=18
+  ad=7290 pd=594 as=0 ps=0
M1467 a_n35820_n12600# s0_not gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1468 a_n31851_n15363# and_a0 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1469 a_n33840_n3285# D vdd w_n33930_n3312# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1470 a_n28026_n9981# a_n29457_n9828# a_n28152_n9981# Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1471 vdd comp_b0 a_n30123_n12375# w_n29898_n12546# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1472 a_n33822_n12447# a3 a_n33822_n12573# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1473 vdd comp_a1 a_n30123_n1953# w_n29898_n2124# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1474 a_n28710_45# a3_not vdd w_n28800_18# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1475 AmoreB_1 a_n28620_n5877# gnd Gnd CMOSN w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
M1476 a_n30123_n3249# comp_b0 a_n30123_n3051# Gnd CMOSN w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1477 a_n29457_n12141# a_n30123_n12177# vdd w_n29547_n11943# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1478 a_n28773_n2844# comp_b0 a_n28377_n2997# Gnd CMOSN w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1479 a_n28773_n2844# x3 vdd w_n28890_n2754# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1480 a_n29565_4599# a_n29286_5148# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1481 and_oper_out2 a_n31851_n14373# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1482 a_n31851_n14499# and_a2 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1483 a1_not comp_a1 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1484 a_n29286_9360# carry2 a_n29286_9234# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1485 and_a3 a_n33822_n12447# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1486 gnd a_n29673_3897# a_n28791_3699# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1487 a_n33822_n14877# D3 vdd w_n33912_n14904# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1488 AequalsB a_n26811_n9819# vdd w_n26433_n9810# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1489 a_n33840_n864# a2 a_n33840_n990# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1490 a_n27954_n765# x3 a_n27954_n891# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1491 a_n33840_n369# D vdd w_n33930_n396# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1492 a_n33840_n1278# D vdd w_n33930_n1305# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1493 vdd comp_a3 a_n30330_n9351# w_n29898_n9288# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1494 comp_b0 a_n30330_n7812# a_n30123_n7380# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1495 a_n29637_4725# a_n29853_5013# vdd w_n29718_4707# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1496 a_n29565_2664# a_n29286_3213# vdd w_n28908_3222# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1497 a_n30123_n6282# a_n30330_n6516# a_n30123_n6084# w_n29898_n6453# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1498 carry3 a_n29637_8820# gnd Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1499 a_n27954_n765# a_n28323_n837# vdd w_n28044_n792# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1500 a_n30312_4959# a_n30483_5832# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1501 a_n28782_n5094# comp_a2 vdd w_n28872_n5121# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1502 a_n28647_n2997# x1 a_n28773_n2997# Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1503 a_n28791_9846# carry2 sum3 Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1504 a_n28710_n4410# b3_not gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1505 a_n30312_9297# adsub_a3 vdd w_n30402_9270# CMOSP w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1506 a_n29637_2790# a_n29853_3078# vdd w_n29718_2772# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1507 x2 a_n30123_n738# vdd w_n29547_n504# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1508 a_n30312_9171# a_n30483_10044# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1509 a_n28782_n765# comp_b2 a_n28683_n891# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1510 D3 a_n35820_n12888# vdd w_n35442_n12879# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1511 a_n30123_n4320# a_n30330_n4554# a_n30123_n4122# w_n29898_n4491# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1512 b2_not comp_b2 gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1513 a_n33822_n11583# b0 a_n33822_n11709# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1514 vdd comp_a1 a_n30330_n6516# w_n29898_n6453# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1515 comp_b1 comp_a1 a_n30123_n10881# w_n29898_n11250# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1516 gnd comp_a3 a_n30123_9# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1517 a_n28620_n5877# x3 vdd w_n28737_n5787# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1518 a_n27072_n5103# AmoreB_2 vdd w_n27576_n5085# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1519 a_n29565_2664# a_n29286_3213# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1520 D a_n34407_n1233# vdd w_n34488_n1134# CMOSP w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1521 vdd adsub_a1 a_n29880_5400# w_n29448_5463# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1522 gnd comp_a0 a_n30123_n3249# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1523 a_n29637_4608# a_n29853_5013# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1524 a_n33822_n12942# D3 vdd w_n33912_n12969# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1525 a_n30123_n936# comp_b2 a_n30123_n738# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1526 gnd comp_a1 a_n30330_n11313# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1527 a_n28620_n1548# x3 vdd w_n28737_n1458# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1528 gnd comp_b1 a_n30330_n2187# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1529 a_n28620_n1701# a1_not gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1530 vdd carry2 a_n28998_9612# w_n28566_9675# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1531 AmoreB_0 a_n28773_n7173# gnd Gnd CMOSN w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
M1532 vdd adsub_a0 a_n29880_3465# w_n29448_3528# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1533 and_oper_out1 a_n31851_n14769# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1534 a_n31851_n14895# and_a1 gnd Gnd CMOSN w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1535 a_n28773_n7173# x2 vdd w_n28890_n7083# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1536 a_n33822_n9135# a1 a_n33822_n9261# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1537 gnd comp_b2 a_n30123_n5265# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1538 adsub_b0 a_n33840_n3816# vdd w_n33462_n3807# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1539 a_n33822_n9666# a0 vdd w_n33912_n9693# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1540 a_n29637_2673# a_n29853_3078# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1541 adsub_b1 a_n33840_n3285# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1542 a_n33822_n15948# D3 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1543 comp_b3 a_n30330_n9351# a_n30123_n8919# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1544 s0_not s0 vdd w_n36243_n12096# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1545 gnd comp_b2 a_n30123_n10062# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1546 AmoreB a_n27072_n5220# vdd w_n27576_n5085# CMOSP w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1547 a_n33822_n14382# b3 vdd w_n33912_n14409# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1548 a_n31851_n15237# and_b0 a_n31851_n15363# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1549 a_n30123_n936# a_n30330_n1170# a_n30123_n738# w_n29898_n1107# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1550 vdd a_n30483_10044# a_n29673_9846# w_n29448_9675# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1551 D1 a_n30690_7515# a_n30483_7947# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1552 a_n28620_n5877# comp_a1 vdd w_n28737_n5787# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1553 a_n35703_n13014# s0 a_n35820_n13014# Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1554 and_b3 a_n33822_n14382# vdd w_n33444_n14373# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1555 a_n29637_6723# a_n29565_6714# a_n29637_6840# w_n29718_6822# CMOSP w=45 l=18
+  ad=1215 pd=144 as=0 ps=0
M1556 and_oper_out3 a_n31851_n13896# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1557 gnd comp_b0 a_n30123_n7578# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1558 a_n28152_n9828# a_n29457_n10845# vdd w_n28260_n9846# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1559 a_n29673_5634# a_n29880_5400# a_n29673_5832# w_n29448_5463# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1560 a_n28620_n1548# comp_b1 vdd w_n28737_n1458# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1561 gnd adsub_a3 a_n29880_9612# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1562 a_n31851_n14373# and_b2 a_n31851_n14499# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1563 a_n33822_n8226# D2 vdd w_n33912_n8253# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1564 adsub_a1 a_n33840_n1278# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1565 a_n33822_n12942# a2 a_n33822_n13068# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1566 s1_not s1 vdd w_n36234_n12420# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1567 a_n33840_n2871# b2 a_n33840_n2997# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1568 a_n33840_n2871# D vdd w_n33930_n2898# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1569 a_n30123_n10062# comp_a2 a_n30123_n9864# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1570 vdd adsub_b3 a_n30690_9612# w_n30258_9675# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1571 vdd comp_a3 a_n30330_n4554# w_n29898_n4491# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1572 a_n29286_9360# a_n29673_10044# vdd w_n29376_9333# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1573 AlessB_2 a_n27954_n765# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1574 a_n27072_n5220# AmoreB_0 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1575 vdd a_n29673_7947# a_n28791_7749# w_n28566_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1576 adsub_a2 a_n33840_n864# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1577 a_n33840_n3285# b1 vdd w_n33930_n3312# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1578 a_n28710_n4284# b3_not vdd w_n28800_n4311# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1579 a_n35820_n12474# s0_not vdd w_n35910_n12501# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1580 gnd carry2 a_n28998_9612# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1581 a_n29637_6723# a_n29565_6714# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1582 comp_a3 comp_b3 a_n30123_207# w_n29898_n162# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1583 b3_not comp_b3 vdd w_n29178_n4194# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1584 a_n29457_n10845# a_n30123_n10881# vdd w_n29547_n10647# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1585 a_n35820_n12888# s0 vdd w_n35910_n12915# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1586 a_n29457_n7344# a_n30123_n7380# vdd w_n29547_n7146# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1587 a_n30483_10044# adsub_a3 a_n29673_10044# w_n29448_9675# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1588 a_n29853_5013# a_n30312_5085# vdd w_n29934_5094# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1589 a_n26982_n774# AlessB_3 a_n27018_n774# w_n27144_n792# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1590 a_n28773_n2844# comp_b0 vdd w_n28890_n2754# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1591 a_n31851_n14373# and_a2 vdd w_n31941_n14400# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1592 a_n28323_n837# a_n28782_n765# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1593 a_n33822_n15003# D3 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1594 a_n29673_3699# a_n29880_3465# a_n29673_3897# w_n29448_3528# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1595 a_n33840_n864# a2 vdd w_n33930_n891# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1596 a_n33822_n11583# b0 vdd w_n33912_n11610# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1597 comp_a1 a_n33822_n9135# vdd w_n33444_n9126# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1598 gnd a_n30483_7947# a_n29673_7749# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1599 comp_b1 a_n30330_n6516# a_n30123_n6084# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1600 a_n33840_n1278# a1 vdd w_n33930_n1305# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1601 a_n33822_n15291# b1 a_n33822_n15417# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1602 a_n29565_6714# a_n29286_7263# vdd w_n28908_7272# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1603 vdd comp_a1 a_n30330_n11313# w_n29898_n11250# CMOSP w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1604 comp_b0 a_n33822_n11583# vdd w_n33444_n11574# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1605 a_n30483_5832# adsub_a1 a_n29673_5832# w_n29448_5463# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1606 comp_b1 a_n33822_n11052# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1607 a_n29286_9234# a_n29673_10044# gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1608 comp_a1 a_n30330_n2187# a_n30123_n1755# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1609 a_n33840_n990# D gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1610 a_n31851_n14769# and_b1 a_n31851_n14895# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1611 a_n28710_n4284# comp_a3 a_n28611_n4410# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1612 vdd D1 a_n30483_7749# w_n30258_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1613 a_n33822_n13356# a1 a_n33822_n13482# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1614 a_n27072_n891# AlessB_0 a_n26892_n774# w_n27144_n792# CMOSP w=45 l=18
+  ad=1215 pd=144 as=0 ps=0
M1615 a_n33822_n13887# a0 vdd w_n33912_n13914# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1616 vdd comp_b2 a_n30123_n10062# w_n29898_n10233# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1617 a_n33822_n10143# b3 a_n33822_n10269# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1618 comp_b3 a_n30330_n4554# a_n30123_n4122# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1619 a_n28773_n2844# x1 vdd w_n28890_n2754# CMOSP w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1620 a_n27072_n774# AlessB_2 vdd w_n27144_n792# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1621 carry3 a_n29637_8820# vdd w_n29718_8919# CMOSP w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1622 a_n28710_45# comp_b3 vdd w_n28800_18# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1623 a_n33840_n3942# D gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1624 and_a0 a_n33822_n13887# vdd w_n33444_n13878# CMOSP w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1625 AmoreB_0 a_n28773_n7173# vdd w_n28890_n7083# CMOSP w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1626 a_n35820_n11565# s1_not a_n35820_n11691# Gnd CMOSN w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1627 and_a1 a_n33822_n13356# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1628 a_n27072_n5220# AmoreB_1 gnd Gnd CMOSN w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1629 comp_b2 comp_a2 a_n30123_n5067# w_n29898_n5436# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1630 a_n29853_5013# a_n30312_5085# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1631 and_oper_out0 a_n31851_n15237# gnd Gnd CMOSN w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1632 a_n30312_9297# a_n30483_10044# vdd w_n30402_9270# CMOSP w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1633 gnd a_n29673_7947# a_n28791_7749# Gnd CMOSN w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1634 a_n28791_7749# a_n28998_7515# sum2 w_n28566_7578# CMOSP w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1635 AlessB_1 a_n28620_n1548# gnd Gnd CMOSN w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
C0 a1 b2 0.82fF
C1 a0 b3 0.82fF
C2 w_n28890_n2754# vdd 11.51fF
C3 w_n33912_n9693# D2 0.93fF
C4 w_n31473_n14364# and_oper_out2 0.19fF
C5 vdd a_n28710_n4284# 0.41fF
C6 D1 sum0 0.99fF
C7 vdd a_n29286_5148# 0.60fF
C8 a_n30483_10044# w_n30258_9675# 1.20fF
C9 adsub_b3 adsub_a2 0.41fF
C10 a_n33840_n3285# b1 0.60fF
C11 vdd a_n29565_2664# 0.60fF
C12 w_n36243_n12096# s0 0.66fF
C13 w_n33912_n12474# vdd 0.28fF
C14 w_n29547_n8685# a_n30123_n8919# 0.66fF
C15 w_n29898_n9288# a_n30123_n9117# 0.72fF
C16 b1 D3 0.13fF
C17 a_n31851_n13896# and_b3 0.60fF
C18 carry2 carry1 0.60fF
C19 a_n28998_3465# sum0 0.99fF
C20 w_n29547_n5850# a_n30123_n6084# 0.66fF
C21 vdd b0 0.27fF
C22 gnd comp_b0 4.26fF
C23 w_n29898_n6453# a_n30123_n6282# 0.72fF
C24 w_n28737_n5787# b1_not 0.63fF
C25 w_n33462_n1800# vdd 1.86fF
C26 a_n29673_5832# a_n28998_5400# 1.08fF
C27 gnd D 5.33fF
C28 w_n28566_7578# a_n29673_7947# 2.98fF
C29 w_n29718_2772# a_n29565_2664# 3.02fF
C30 w_n33912_n8253# D2 0.93fF
C31 x3 a_n27954_n5094# 1.21fF
C32 a_n28998_9612# carry2 2.85fF
C33 gnd a_n29853_9225# 0.60fF
C34 x3 comp_b1 0.04fF
C35 b1 a_n33822_n15291# 0.60fF
C36 w_n31941_n15264# a_n31851_n15237# 0.42fF
C37 w_n33912_n11610# vdd 0.28fF
C38 w_n29547_n1521# x1 0.19fF
C39 w_n33912_n9162# a1 0.93fF
C40 and_a2 and_b2 0.87fF
C41 w_n33444_n8217# comp_a3 0.19fF
C42 D1 gnd 8.91fF
C43 w_n29205_n675# vdd 1.92fF
C44 w_n29448_7578# a_n29673_7947# 1.20fF
C45 a_n30330_n2187# comp_a1 1.73fF
C46 w_n29547_n2817# x0 0.19fF
C47 w_n29934_3159# a_n30312_3150# 2.17fF
C48 w_n31941_n13923# and_b3 0.93fF
C49 D1 a_n30690_3465# 1.03fF
C50 vdd a_n29673_5832# 1.21fF
C51 vdd s0 0.60fF
C52 AlessB_3 a_n27072_n891# 1.04fF
C53 comp_a1 comp_a0 0.35fF
C54 vdd and_a0 0.77fF
C55 comp_b1 a_n30330_n11313# 0.99fF
C56 comp_b2 a_n30123_n5067# 1.27fF
C57 gnd a_n28998_3465# 0.60fF
C58 w_n35442_n11556# a_n35820_n11565# 2.17fF
C59 w_n33912_n10665# vdd 0.28fF
C60 a_n30330_n5499# a_n30123_n5067# 0.99fF
C61 comp_b2 a_n30123_n9864# 1.27fF
C62 w_n28890_n7083# AmoreB_0 0.19fF
C63 w_n33462_n360# vdd 1.86fF
C64 a_n30330_n10296# a_n30123_n9864# 0.99fF
C65 vdd a_n35820_n12474# 0.60fF
C66 a3 D3 0.04fF
C67 w_n28737_n1458# AlessB_1 0.19fF
C68 vdd a_n30123_n738# 1.04fF
C69 comp_a2 x2 0.92fF
C70 adsub_b1 adsub_a0 0.41fF
C71 gnd comp_b2 5.33fF
C72 vdd comp_a2 1.86fF
C73 b2 a_n33822_n14877# 0.60fF
C74 gnd a_n30330_n5499# 0.60fF
C75 w_n33444_n10134# vdd 1.86fF
C76 w_n29898_n10233# comp_a2 1.86fF
C77 gnd a_n30330_n10296# 0.60fF
C78 x3 a_n28620_n1548# 1.67fF
C79 b1 b0 0.95fF
C80 w_n33912_n8748# a2 0.93fF
C81 gnd b3 3.49fF
C82 w_n28800_n4311# comp_a3 0.93fF
C83 vdd a_n31851_n14769# 0.41fF
C84 w_n30402_3123# vdd 0.28fF
C85 comp_b0 a_n30123_n3051# 0.99fF
C86 vdd a_n29565_6714# 0.60fF
C87 a_n30690_7515# adsub_b2 1.00fF
C88 w_n29448_3528# adsub_a0 1.86fF
C89 vdd a_n33822_n9666# 0.60fF
C90 w_n28566_7578# sum2 1.20fF
C91 a_n28998_5400# sum1 0.99fF
C92 comp_b1 a_n30123_n1953# 1.98fF
C93 vdd a_n33822_n12942# 0.60fF
C94 w_n33444_n14868# and_b2 0.19fF
C95 a_n30330_n225# a_n30123_207# 0.99fF
C96 w_n33444_n10134# a_n33822_n10143# 2.17fF
C97 w_n33444_n8712# vdd 1.86fF
C98 gnd a_n30330_n9351# 0.60fF
C99 w_n29898_n12546# comp_a0 1.86fF
C100 w_n33930_n2403# a_n33840_n2376# 0.42fF
C101 w_n28044_n5121# a_n28323_n5166# 0.93fF
C102 w_n27576_n5085# AmoreB_2 0.99fF
C103 gnd comp_a3 5.43fF
C104 w_n30402_5058# vdd 0.28fF
C105 x3 a_n28620_n5877# 1.67fF
C106 a_n29565_6714# a_n29637_6723# 1.62fF
C107 a_n30330_n9351# a_n30123_n8919# 0.99fF
C108 w_n28872_n792# a_n28782_n765# 0.42fF
C109 x2 a_n28494_n6030# 0.06fF
C110 w_n28737_n5787# x3 0.81fF
C111 comp_a3 a_n30123_n8919# 0.99fF
C112 b3 a_n33822_n14382# 0.60fF
C113 a_n29457_n10845# a_n28152_n9828# 0.80fF
C114 a2 D3 0.10fF
C115 w_n29547_n5850# vdd 1.95fF
C116 comp_b1 a_n30123_n6282# 1.98fF
C117 gnd a_n29853_3078# 0.60fF
C118 w_n30402_7173# vdd 0.28fF
C119 w_n33912_n12474# a3 0.93fF
C120 adsub_a0 a_n29673_3699# 3.02fF
C121 w_n31941_n13923# and_a3 0.93fF
C122 a3 b0 0.82fF
C123 a_n30483_5832# a_n29673_5634# 1.98fF
C124 w_n33912_n15318# vdd 0.28fF
C125 vdd a_n33822_n12447# 0.60fF
C126 w_n29268_n7146# comp_b0 0.66fF
C127 w_n29547_n4833# x2 0.19fF
C128 comp_b0 a_n30123_n7578# 1.98fF
C129 s1_not a_n35820_n11691# 0.06fF
C130 w_n29547_n4833# vdd 2.02fF
C131 w_n29718_6822# a_n29565_6714# 3.02fF
C132 comp_b1 a_n28620_n1701# 0.10fF
C133 vdd a_n28782_n5094# 1.02fF
C134 comp_b3 a_n28710_45# 0.60fF
C135 w_n28566_3528# D1 1.95fF
C136 vdd w_n28908_9369# 1.86fF
C137 vdd a_n29457_n9828# 0.80fF
C138 comp_a2 comp_a1 1.33fF
C139 a_n30690_9612# a_n30483_10044# 0.99fF
C140 gnd x3 1.85fF
C141 w_n33912_n14409# vdd 0.28fF
C142 w_n29898_n3420# a_n30123_n3051# 1.20fF
C143 w_n33912_n13914# a_n33822_n13887# 0.42fF
C144 s1_not a_n35820_n12159# 0.06fF
C145 w_n33444_n13878# and_a0 0.19fF
C146 w_n28566_3528# a_n28998_3465# 1.29fF
C147 w_n33462_n3807# vdd 1.86fF
C148 w_n29934_7209# a_n30312_7200# 2.17fF
C149 w_n31473_n14760# a_n31851_n14769# 2.17fF
C150 w_n33444_n14868# a_n33822_n14877# 2.17fF
C151 w_n29898_n162# a_n30123_207# 1.20fF
C152 comp_b3 comp_a0 0.68fF
C153 adsub_b0 a_n30483_3897# 0.99fF
C154 w_n33462_n2862# a_n33840_n2871# 2.17fF
C155 w_n28737_n5787# AmoreB_1 0.19fF
C156 w_n33444_n13347# vdd 1.86fF
C157 a_n29286_9360# w_n29376_9333# 0.42fF
C158 gnd adsub_b1 1.72fF
C159 gnd a_n30330_n11313# 0.60fF
C160 w_n33462_n2862# vdd 1.86fF
C161 w_n28044_n792# a_n27954_n765# 0.42fF
C162 a2 b0 0.82fF
C163 comp_b2 comp_b0 1.66fF
C164 w_n29376_7236# carry1 0.93fF
C165 w_n29178_135# comp_a3 0.66fF
C166 D1 a_n28998_3465# 2.85fF
C167 a0 D2 0.12fF
C168 a_n29673_10044# a_n28791_9846# 1.98fF
C169 w_n33912_n15318# b1 0.93fF
C170 vdd a1 0.27fF
C171 D b3 0.09fF
C172 w_n35910_n12501# vdd 0.28fF
C173 vdd and_b2 1.80fF
C174 w_n29898_n9288# a_n30123_n8919# 1.20fF
C175 a_n28791_9846# w_n28566_9675# 0.72fF
C176 w_n30258_3528# adsub_b0 1.86fF
C177 gnd a_n29853_7128# 0.60fF
C178 adsub_a0 a_n30312_3150# 1.81fF
C179 w_n29898_n3420# comp_b0 1.86fF
C180 w_n28737_n1458# x2 0.84fF
C181 w_n29898_n6453# a_n30123_n6084# 1.20fF
C182 x3 a_n27954_n765# 1.21fF
C183 w_n28737_n1458# vdd 11.51fF
C184 vdd a_n33840_n3816# 0.60fF
C185 w_n29898_n11250# comp_b1 2.98fF
C186 x1 a_n28773_n7173# 1.58fF
C187 w_n33912_n8253# a_n33822_n8226# 0.42fF
C188 x3 a_n28323_n5166# 0.06fF
C189 D1 w_n30258_9675# 2.98fF
C190 w_n28404_n5085# a_n28782_n5094# 2.17fF
C191 w_n29205_n5004# b2_not 0.19fF
C192 comp_a3 comp_b0 0.48fF
C193 w_n33444_n11574# vdd 1.86fF
C194 gnd AmoreB_1 1.07fF
C195 a_n29673_10044# w_n29376_9333# 0.93fF
C196 w_n29376_5121# a_n29286_5148# 0.42fF
C197 w_n29547_n504# x2 0.19fF
C198 w_n29547_n504# vdd 2.02fF
C199 a_n30690_9612# gnd 0.60fF
C200 w_n30402_7173# adsub_b2 0.05fF
C201 comp_b0 a_n28377_n2997# 0.06fF
C202 w_n30258_7578# D1 2.98fF
C203 w_n31941_n13923# a_n31851_n13896# 0.42fF
C204 a_n29880_7515# adsub_a2 1.03fF
C205 w_n27144_n792# a_n27072_n891# 0.96fF
C206 w_n29547_n10647# a_n30123_n10881# 0.66fF
C207 w_n29898_n11250# a_n30123_n11079# 0.72fF
C208 vdd a_n33822_n13887# 0.60fF
C209 w_n33444_n10629# vdd 1.86fF
C210 comp_b2 a_n30330_n5499# 1.73fF
C211 w_n29214_n1521# a1_not 0.19fF
C212 w_n33912_n13383# D3 0.93fF
C213 w_n28566_5463# a_n28791_5634# 0.72fF
C214 a_n30483_3897# adsub_a0 1.55fF
C215 comp_b2 a_n30330_n10296# 1.06fF
C216 a_n35820_n12474# s1 0.60fF
C217 w_n28800_18# vdd 0.28fF
C218 and_a0 and_b1 0.54fF
C219 gnd adsub_a1 2.41fF
C220 a3 a_n33822_n12447# 0.60fF
C221 b0 a_n33822_n11583# 0.60fF
C222 a1 b1 0.82fF
C223 a0 b2 0.82fF
C224 comp_a2 a_n30123_n936# 1.98fF
C225 a2 a_n33822_n12942# 0.60fF
C226 w_n33912_n9693# vdd 0.28fF
C227 w_n33912_n12474# D3 0.93fF
C228 w_n29376_5121# a_n29673_5832# 0.93fF
C229 x3 comp_b0 0.41fF
C230 vdd a_n33822_n14877# 0.60fF
C231 w_n29934_3159# vdd 1.86fF
C232 a_n30330_n11313# a_n30123_n10881# 0.99fF
C233 w_n33462_n360# adsub_a3 0.19fF
C234 b0 D3 0.06fF
C235 comp_b3 comp_a2 1.33fF
C236 w_n34488_n1134# D 0.14fF
C237 w_n33912_n11610# a_n33822_n11583# 0.42fF
C238 x2 x1 0.27fF
C239 comp_a3 comp_b2 0.34fF
C240 comp_b1 a_n30285_n7686# 0.06fF
C241 w_n33912_n13383# a_n33822_n13356# 0.42fF
C242 w_n33444_n13347# and_a1 0.19fF
C243 vdd x1 1.23fF
C244 w_n33444_n10134# comp_b3 0.19fF
C245 w_n29448_3528# a_n29880_3465# 1.29fF
C246 gnd D2 4.84fF
C247 adsub_a1 a_n30312_5085# 1.81fF
C248 comp_b1 a_n30123_n1755# 0.99fF
C249 w_n29898_n4491# a_n30123_n4320# 0.72fF
C250 w_n29547_n3888# a_n30123_n4122# 0.66fF
C251 a_n31851_n14769# and_b1 0.60fF
C252 w_n33912_n8253# vdd 0.28fF
C253 w_n33462_n2862# adsub_b2 0.19fF
C254 vdd a_n29286_9360# 0.60fF
C255 w_n27576_n5085# a_n27954_n5094# 2.17fF
C256 w_n33462_n2367# a_n33840_n2376# 2.17fF
C257 w_n34488_n1134# D1 0.80fF
C258 w_n29934_5094# vdd 1.86fF
C259 w_n36234_n12420# s1_not 0.19fF
C260 gnd a_n30330_n225# 0.60fF
C261 w_n33912_n11079# a_n33822_n11052# 0.42fF
C262 and_a1 and_b2 0.54fF
C263 w_n33930_n3843# b0 0.93fF
C264 a_n29880_9612# adsub_a3 1.03fF
C265 w_n28044_n5121# x3 2.64fF
C266 w_n30402_7173# adsub_a2 0.93fF
C267 w_n33930_n891# a_n33840_n864# 0.42fF
C268 w_n31941_n15264# and_a0 0.93fF
C269 D1 a_n30483_3699# 1.98fF
C270 w_n29898_n6453# vdd 0.48fF
C271 w_n33912_n9162# a_n33822_n9135# 0.42fF
C272 comp_b1 a_n30123_n6084# 1.27fF
C273 vdd a_n33822_n11052# 0.60fF
C274 vdd D0 1.04fF
C275 a3 a1 0.82fF
C276 w_n35910_n11592# s1_not 0.93fF
C277 w_n29934_7209# vdd 1.86fF
C278 w_n28800_18# a3_not 0.93fF
C279 D1 adsub_b1 0.11fF
C280 w_n33462_n1269# adsub_a1 0.19fF
C281 adsub_a0 a_n29673_3897# 2.03fF
C282 w_n33444_n15282# vdd 1.86fF
C283 a_n30483_5832# a_n29673_5832# 0.99fF
C284 x3 comp_b2 0.04fF
C285 w_n28890_n7083# x1 0.74fF
C286 AmoreB_1 a_n27072_n5220# 1.06fF
C287 gnd carry0 1.21fF
C288 vdd a_n28782_n765# 1.02fF
C289 comp_b0 a_n30123_n7380# 1.27fF
C290 w_n29898_n5436# vdd 0.48fF
C291 vdd a_n29673_10044# 1.21fF
C292 w_n27576_n5085# AmoreB_3 2.24fF
C293 vdd w_n28566_9675# 0.48fF
C294 w_n28737_n1458# temp_less 0.63fF
C295 and_a2 and_b3 0.54fF
C296 gnd b2 3.55fF
C297 w_n31473_n14364# vdd 1.14fF
C298 w_n29547_n9630# a_n30123_n9864# 0.66fF
C299 vdd a_n30123_207# 1.04fF
C300 w_n29898_n10233# a_n30123_n10062# 0.72fF
C301 comp_b0 a_n28773_n2844# 0.80fF
C302 w_n33444_n13878# a_n33822_n13887# 2.17fF
C303 comp_a2 comp_a0 15.88fF
C304 adsub_b2 a_n30483_7749# 1.98fF
C305 w_n29268_n2817# vdd 1.62fF
C306 adsub_a3 a_n29673_9846# 2.83fF
C307 s0_not s1_not 4.35fF
C308 comp_a1 x1 1.23fF
C309 w_n33912_n11610# b0 0.93fF
C310 vdd adsub_b0 0.76fF
C311 gnd a_n30483_3897# 0.74fF
C312 comp_a3 x3 0.99fF
C313 comp_b3 a_n30123_9# 1.98fF
C314 w_n29898_n2124# comp_b1 1.86fF
C315 carry2 a_n29286_9360# 1.81fF
C316 a_n30690_3465# a_n30483_3897# 0.99fF
C317 a_n30690_9612# D1 1.06fF
C318 a2 a1 0.82fF
C319 w_n33912_n12969# vdd 0.28fF
C320 w_n29547_n8685# a_n29457_n8883# 0.19fF
C321 a_n29853_9225# w_n29718_8919# 0.80fF
C322 a_n29565_8811# w_n28908_9369# 0.19fF
C323 gnd a_n30690_5400# 0.60fF
C324 b1 a_n33822_n11052# 0.60fF
C325 w_n28044_n792# a_n28323_n837# 0.93fF
C326 w_n33930_n2403# vdd 0.28fF
C327 w_n27576_n756# AlessB_2 0.19fF
C328 w_n33912_n13914# a0 0.93fF
C329 gnd and_a2 0.60fF
C330 vdd a_n30123_n4122# 1.04fF
C331 a_n28998_7515# carry1 2.85fF
C332 comp_a1 a_n28620_n6030# 0.10fF
C333 w_n35910_n12501# s1 0.93fF
C334 w_n30402_5058# a_n30483_5832# 0.93fF
C335 vdd a_n33840_n1278# 0.60fF
C336 w_n28044_n792# x3 2.64fF
C337 vdd a_n29286_3213# 0.60fF
C338 vdd a_n31851_n14373# 0.41fF
C339 w_n36234_n12420# vdd 2.50fF
C340 w_n29898_n6453# comp_a1 1.86fF
C341 w_n29898_n9288# a_n30330_n9351# 1.29fF
C342 w_n33912_n15318# D3 0.93fF
C343 a_n29673_3897# sum0 1.55fF
C344 comp_b3 a_n30123_n4320# 1.98fF
C345 D1 adsub_a1 0.12fF
C346 w_n33444_n12933# and_a2 0.19fF
C347 w_n30258_3528# a_n30690_3465# 1.29fF
C348 w_n29898_n9288# comp_a3 1.86fF
C349 w_n29898_n6453# a_n30330_n6516# 1.29fF
C350 x3 a_n28323_n837# 0.06fF
C351 w_n33930_n1305# vdd 0.28fF
C352 vdd AlessB_3 0.60fF
C353 w_n33930_n3312# D 0.93fF
C354 w_n33444_n8217# a_n33822_n8226# 2.17fF
C355 a_n30690_9612# w_n30258_9675# 1.29fF
C356 gnd AlessB_1 1.07fF
C357 w_n33912_n8253# a3 0.93fF
C358 gnd a_n30285_n7686# 1.49fF
C359 a_n29673_10044# carry2 0.09fF
C360 vdd a_n27954_n5094# 0.60fF
C361 w_n33912_n15318# a_n33822_n15291# 0.42fF
C362 w_n35910_n11592# vdd 0.28fF
C363 w_n36243_n12096# s0_not 0.19fF
C364 x2 comp_b1 0.04fF
C365 carry2 w_n28566_9675# 1.95fF
C366 vdd comp_b1 2.71fF
C367 w_n33912_n14409# D3 0.93fF
C368 w_n28908_5157# a_n29565_4599# 0.19fF
C369 w_n29547_n11943# a_n30123_n12177# 0.66fF
C370 w_n29718_4707# a_n29853_5013# 0.80fF
C371 w_n29898_n12546# a_n30123_n12375# 0.72fF
C372 w_n35910_n12915# a_n35820_n12888# 0.42fF
C373 adsub_b3 a_n30483_9846# 1.98fF
C374 w_n29898_n1107# vdd 0.48fF
C375 w_n29205_n675# comp_a2 0.66fF
C376 w_n31473_n13887# a_n31851_n13896# 2.17fF
C377 w_n29898_n11250# a_n30123_n10881# 1.20fF
C378 a3 D0 0.06fF
C379 w_n29547_441# x3 0.19fF
C380 gnd a_n29673_3897# 1.02fF
C381 vdd adsub_a0 1.81fF
C382 w_n26901_n9846# vdd 0.28fF
C383 gnd a_n29457_n12141# 0.80fF
C384 vdd a_n30483_7947# 0.60fF
C385 a_n30483_3897# a_n29880_3465# 1.60fF
C386 a_n30330_n3483# comp_a0 1.73fF
C387 w_n28332_54# vdd 1.14fF
C388 gnd and_b0 1.20fF
C389 gnd a_n29880_5400# 0.60fF
C390 w_n27144_n792# AlessB_1 0.99fF
C391 comp_a2 a_n30123_n738# 1.27fF
C392 a_n33840_n2376# b3 0.60fF
C393 vdd s0_not 0.73fF
C394 gnd s1_not 1.35fF
C395 D1 a_n34407_n1233# 0.60fF
C396 vdd AmoreB_3 0.60fF
C397 w_n28800_18# comp_b3 0.93fF
C398 a1 D3 0.10fF
C399 w_n33444_n9657# vdd 1.86fF
C400 w_n33912_n12474# a_n33822_n12447# 0.42fF
C401 w_n29898_n12546# a_n30330_n12609# 1.29fF
C402 b3 D2 0.12fF
C403 vdd a0 0.27fF
C404 w_n28566_5463# carry0 1.95fF
C405 D b2 0.12fF
C406 w_n28908_3222# vdd 1.86fF
C407 w_n33444_n11574# a_n33822_n11583# 2.17fF
C408 x2 a_n28620_n1548# 1.16fF
C409 w_n33930_n891# D 0.93fF
C410 w_n35910_n12060# a_n35820_n12033# 0.42fF
C411 D1 carry0 0.46fF
C412 w_n33444_n13347# a_n33822_n13356# 2.17fF
C413 vdd a_n29286_7263# 0.60fF
C414 vdd a_n33822_n9135# 0.60fF
C415 a_n30483_10044# vdd 0.60fF
C416 a_n29673_5832# sum1 1.55fF
C417 w_n29898_n4491# a_n30123_n4122# 1.20fF
C418 vdd a_n30123_n12177# 1.04fF
C419 w_n31941_n14400# and_b2 0.93fF
C420 w_n33444_n8217# vdd 1.86fF
C421 w_n33444_n8712# comp_a2 0.19fF
C422 comp_b3 x1 0.41fF
C423 carry2 sum3 0.99fF
C424 a2 D0 0.06fF
C425 w_n28908_5157# vdd 1.86fF
C426 w_n33444_n11043# a_n33822_n11052# 2.17fF
C427 a1 a_n33822_n13356# 0.60fF
C428 x3 a_n28773_n2844# 1.16fF
C429 w_n33930_n3843# a_n33840_n3816# 0.42fF
C430 w_n28404_n756# a_n28782_n765# 2.17fF
C431 w_n29205_n675# a2_not 0.19fF
C432 x2 a_n28620_n5877# 1.16fF
C433 w_n28872_n792# comp_b2 0.93fF
C434 w_n33912_n13383# a1 0.93fF
C435 comp_a1 comp_b1 0.80fF
C436 w_n33462_n855# a_n33840_n864# 2.17fF
C437 a_n29457_n9828# a_n28152_n9828# 0.80fF
C438 adsub_a2 a_n29673_7749# 2.83fF
C439 D1 a_n30483_3897# 0.99fF
C440 a_n30330_n225# comp_a3 1.80fF
C441 w_n28737_n5787# x2 0.84fF
C442 w_n28890_n2754# AlessB_0 0.19fF
C443 w_n33444_n9126# a_n33822_n9135# 2.17fF
C444 w_n28737_n5787# vdd 11.51fF
C445 comp_b1 a_n30330_n6516# 1.73fF
C446 vdd a_n33840_n864# 0.60fF
C447 vdd and_b3 1.06fF
C448 w_n35442_n12465# D2 0.19fF
C449 w_n28800_18# a_n28710_45# 0.42fF
C450 w_n28908_7272# vdd 1.86fF
C451 D1 a_n30690_5400# 1.06fF
C452 vdd a_n29673_7947# 1.21fF
C453 a_n29880_3465# a_n29673_3897# 0.99fF
C454 w_n31473_n15228# vdd 1.14fF
C455 w_n28260_n9846# temp 0.63fF
C456 gnd a_n28998_5400# 0.60fF
C457 w_n29898_n7749# comp_b0 2.98fF
C458 w_n28800_n4311# vdd 0.28fF
C459 comp_b0 a_n30285_n7686# 0.75fF
C460 a0 b1 0.82fF
C461 a1 b0 0.82fF
C462 b3 b2 1.08fF
C463 comp_a1 a_n30123_n11079# 1.98fF
C464 w_n30258_3528# D1 2.98fF
C465 w_n33444_n15282# and_b1 0.19fF
C466 vdd a_n30123_n5067# 1.04fF
C467 comp_a2 a_n28782_n5094# 0.60fF
C468 vdd w_n29448_9675# 0.48fF
C469 w_n29898_n7749# a_n30123_n7578# 0.72fF
C470 w_n28890_n7083# b0_not 0.63fF
C471 w_n29547_n7146# a_n30123_n7380# 0.66fF
C472 a_n33840_n3816# b0 0.60fF
C473 a_n30285_n7686# a_n30123_n7578# 1.98fF
C474 vdd a_n30123_n9864# 1.04fF
C475 w_n27576_n5085# a_n27072_n5220# 0.96fF
C476 w_n33444_n14373# vdd 1.86fF
C477 w_n28260_n9846# a_n29457_n8883# 0.63fF
C478 vdd a_n33840_n369# 0.60fF
C479 adsub_b2 adsub_a0 0.41fF
C480 w_n29898_n10233# a_n30123_n9864# 1.20fF
C481 carry3 w_n29718_8919# 0.14fF
C482 w_n33912_n12969# a2 0.93fF
C483 w_n28890_n2754# a0_not 0.63fF
C484 w_n28566_3528# a_n29673_3897# 2.98fF
C485 adsub_b2 a_n30483_7947# 1.16fF
C486 w_n29448_3528# a_n29673_3699# 0.72fF
C487 w_n29547_n2817# vdd 1.95fF
C488 gnd x2 1.31fF
C489 a_n35820_n11565# s1_not 0.60fF
C490 gnd vdd 14.95fF
C491 adsub_a3 a_n29673_10044# 1.84fF
C492 carry0 a_n28791_5634# 1.98fF
C493 w_n30258_5463# D1 2.98fF
C494 comp_b3 a_n30123_207# 0.99fF
C495 a_n29673_7947# a_n28791_7749# 1.98fF
C496 a_n30483_10044# w_n30402_9270# 0.93fF
C497 vdd a_n30123_n8919# 1.04fF
C498 x1 comp_a0 0.41fF
C499 w_n33444_n12933# vdd 1.86fF
C500 and_a0 and_b2 0.54fF
C501 comp_a0 a_n30123_n12375# 1.98fF
C502 w_n27576_n756# a_n27954_n765# 2.17fF
C503 w_n33462_n2367# vdd 1.86fF
C504 comp_b3 a_n30123_n9117# 0.99fF
C505 w_n34488_n1134# a_n34407_n1233# 0.96fF
C506 w_n26433_n9810# AequalsB 0.19fF
C507 vdd a_n30312_5085# 0.60fF
C508 adsub_b3 adsub_a0 0.41fF
C509 D1 a_n29673_3897# 0.09fF
C510 w_n29898_n162# comp_a3 2.98fF
C511 comp_a1 a_n28620_n5877# 0.80fF
C512 w_n36234_n12420# s1 0.66fF
C513 w_n29448_5463# adsub_a1 1.86fF
C514 w_n35910_n12501# a_n35820_n12474# 0.42fF
C515 comp_b2 a_n30285_n7686# 0.27fF
C516 a3 a0 0.82fF
C517 vdd a_n33822_n14382# 0.60fF
C518 w_n33444_n12438# vdd 1.86fF
C519 w_n28737_n5787# comp_a1 0.63fF
C520 w_n28890_n2754# x1 0.74fF
C521 comp_b3 a_n30123_n4122# 1.27fF
C522 a_n29673_3897# a_n28998_3465# 1.08fF
C523 w_n27144_n792# vdd 3.84fF
C524 w_n26901_n9846# k 0.93fF
C525 w_n33444_n11043# comp_b1 0.19fF
C526 vdd and_a3 0.62fF
C527 w_n29376_3186# a_n29286_3213# 0.42fF
C528 s1_not a_n35820_n12033# 0.60fF
C529 vdd a_n27954_n765# 0.60fF
C530 gnd a_n30330_n7812# 0.60fF
C531 w_n33930_n1836# a0 0.93fF
C532 a_n29673_10044# a_n28998_9612# 1.08fF
C533 w_n33444_n15282# a_n33822_n15291# 2.17fF
C534 w_n31473_n15228# a_n31851_n15237# 2.17fF
C535 temp_less a_n28620_n1548# 0.80fF
C536 w_n35442_n11556# vdd 1.86fF
C537 a_n28998_9612# w_n28566_9675# 1.29fF
C538 w_n29547_n7146# a_n29457_n7344# 0.19fF
C539 and_a1 and_b3 0.54fF
C540 w_n35442_n12879# a_n35820_n12888# 2.17fF
C541 w_n29898_n12546# a_n30123_n12177# 1.20fF
C542 w_n29898_n1107# a_n30123_n936# 0.72fF
C543 w_n29547_n504# a_n30123_n738# 0.66fF
C544 gnd b1 3.57fF
C545 adsub_b3 a_n30483_10044# 1.16fF
C546 w_n33462_n1269# vdd 1.86fF
C547 comp_a3 a_n30285_n7686# 0.01fF
C548 vdd a_n30123_n3051# 1.04fF
C549 a_n30483_7947# adsub_a2 1.43fF
C550 w_n28566_3528# a_n28791_3699# 0.72fF
C551 comp_b3 comp_b1 1.47fF
C552 gnd carry2 1.21fF
C553 w_n29898_n11250# a_n30330_n11313# 1.29fF
C554 w_n31473_n14760# and_oper_out1 0.19fF
C555 w_n26433_n9810# vdd 1.14fF
C556 gnd comp_a1 5.67fF
C557 gnd a_n29457_n10845# 0.80fF
C558 w_n33912_n12969# D3 0.93fF
C559 b2 a_n33822_n10638# 0.60fF
C560 a2 a0 0.82fF
C561 gnd a_n30330_n6516# 0.60fF
C562 w_n29178_135# vdd 1.86fF
C563 w_n29268_n2817# comp_a0 0.66fF
C564 vdd a_n30123_n10881# 1.04fF
C565 vdd a_n35820_n11565# 0.60fF
C566 D0 b0 0.10fF
C567 w_n28800_n4311# b3_not 0.93fF
C568 gnd and_a1 0.60fF
C569 D1 a_n28791_3699# 1.98fF
C570 w_n29547_n8685# vdd 2.02fF
C571 gnd adsub_b2 1.72fF
C572 w_n28566_5463# a_n28998_5400# 1.29fF
C573 vdd a_n33840_n1809# 0.60fF
C574 temp_more a_n28620_n5877# 0.80fF
C575 a_n30690_5400# adsub_b1 1.00fF
C576 w_n28566_3528# vdd 0.48fF
C577 a_n33840_n369# a3 0.60fF
C578 w_n29214_n5850# comp_b1 0.66fF
C579 w_n29448_3528# a_n30483_3897# 2.98fF
C580 comp_a2 x1 0.04fF
C581 w_n30258_3528# a_n30483_3699# 0.72fF
C582 comp_b0 x2 0.41fF
C583 w_n28737_n5787# temp_more 0.63fF
C584 vdd comp_b0 2.34fF
C585 gnd a3 2.62fF
C586 w_n29898_n4491# a_n30330_n4554# 1.29fF
C587 w_n31941_n14400# a_n31851_n14373# 0.42fF
C588 w_n33912_n9693# a_n33822_n9666# 0.42fF
C589 w_n29268_n7146# vdd 1.62fF
C590 a_n28998_9612# sum3 0.99fF
C591 a_n29565_4599# a_n29637_4608# 1.62fF
C592 w_n28404_n5085# a_n28323_n5166# 0.19fF
C593 a2 a_n33840_n864# 0.60fF
C594 w_n28566_5463# vdd 0.48fF
C595 w_n33462_n3807# a_n33840_n3816# 2.17fF
C596 a_n30483_10044# adsub_a3 1.43fF
C597 adsub_b3 gnd 1.72fF
C598 D1 vdd 2.17fF
C599 a_n30330_n2187# comp_b1 2.31fF
C600 adsub_a2 a_n29673_7947# 1.84fF
C601 w_n28044_n5121# vdd 0.28fF
C602 vdd a_n35820_n12033# 0.60fF
C603 w_n30258_5463# adsub_b1 1.86fF
C604 w_n33912_n14904# b2 0.93fF
C605 comp_b1 comp_a0 0.40fF
C606 vdd a_n31851_n13896# 0.41fF
C607 w_n28332_54# a_n28710_45# 2.17fF
C608 w_n29178_135# a3_not 0.19fF
C609 w_n28566_7578# vdd 0.48fF
C610 AlessB_1 a_n27072_n891# 1.06fF
C611 a_n30483_3897# a_n29673_3699# 1.98fF
C612 w_n33462_n2367# adsub_b3 0.19fF
C613 comp_a0 a_n30123_n3249# 1.98fF
C614 w_n31941_n14796# vdd 0.28fF
C615 w_n29547_n3888# x3 0.23fF
C616 w_n26901_n9846# a_n26811_n9819# 0.42fF
C617 w_n28260_n9846# a_n29457_n12141# 0.63fF
C618 w_n29547_n5850# x1 0.19fF
C619 comp_b0 a_n30330_n7812# 1.73fF
C620 w_n28332_n4275# vdd 1.14fF
C621 comp_b2 x2 0.90fF
C622 w_n29898_n5436# comp_a2 1.86fF
C623 gnd a2 2.48fF
C624 vdd comp_b2 1.86fF
C625 w_n29376_7236# a_n29286_7263# 0.42fF
C626 comp_a1 a_n30123_n10881# 0.99fF
C627 w_n33930_n396# a_n33840_n369# 0.42fF
C628 w_n29448_7578# vdd 0.48fF
C629 w_n29898_n7749# a_n30123_n7380# 1.20fF
C630 carry1 a_n29286_7263# 1.81fF
C631 a0 D3 0.10fF
C632 comp_a2 a_n30123_n5265# 1.98fF
C633 vdd w_n30258_9675# 0.48fF
C634 w_n29898_n10233# comp_b2 2.98fF
C635 gnd adsub_a2 2.13fF
C636 b2 D2 0.12fF
C637 comp_a2 a_n30123_n10062# 1.98fF
C638 a_n30285_n7686# a_n30123_n7380# 0.99fF
C639 vdd b3 0.27fF
C640 D b1 0.09fF
C641 w_n31941_n13923# vdd 0.28fF
C642 w_n29898_n10233# a_n30330_n10296# 1.29fF
C643 x2 a_n28494_n1701# 0.06fF
C644 gnd s1 2.01fF
C645 a_n29637_8820# w_n29718_8919# 0.96fF
C646 a_n30690_7515# a_n30483_7947# 0.99fF
C647 w_n29448_3528# a_n29673_3897# 1.20fF
C648 w_n29898_n3420# vdd 0.48fF
C649 a_n29880_9612# a_n29673_10044# 0.99fF
C650 x3 a_n28773_n7173# 1.16fF
C651 w_n33444_n9657# comp_a0 0.19fF
C652 w_n28566_7578# a_n28791_7749# 0.72fF
C653 w_n30258_7578# vdd 0.48fF
C654 adsub_a3 w_n29448_9675# 1.86fF
C655 comp_b0 comp_a1 0.16fF
C656 w_n27576_n5085# AmoreB_1 0.99fF
C657 b3 a_n33822_n10143# 0.60fF
C658 D1 b1 0.58fF
C659 comp_a3 x2 0.04fF
C660 gnd and_b1 0.60fF
C661 vdd comp_a3 2.20fF
C662 w_n35910_n12915# vdd 0.28fF
C663 gnd comp_b3 5.33fF
C664 a_n29286_9360# w_n28908_9369# 2.17fF
C665 w_n33462_n3276# adsub_b1 0.19fF
C666 comp_a0 a_n30123_n12177# 0.99fF
C667 w_n29214_n1521# vdd 1.29fF
C668 adsub_a3 gnd 1.67fF
C669 comp_b3 a_n30123_n8919# 1.27fF
C670 w_n29376_7236# a_n29673_7947# 0.93fF
C671 w_n33462_n1800# adsub_a0 0.19fF
C672 a_n26811_n9819# equals_d 0.60fF
C673 w_n29898_n162# a_n30330_n225# 1.29fF
C674 w_n33912_n9162# D2 0.93fF
C675 a_n29673_7947# carry1 0.09fF
C676 w_n29448_5463# a_n29880_5400# 1.29fF
C677 w_n35442_n12465# vdd 1.86fF
C678 D1 a_n30483_5634# 1.98fF
C679 w_n33912_n12969# a_n33822_n12942# 0.42fF
C680 comp_b3 a_n30330_n4554# 1.73fF
C681 w_n29718_4707# a_n29637_4608# 0.96fF
C682 w_n28044_n792# vdd 0.28fF
C683 w_n33930_n2898# D 0.93fF
C684 D a3 0.04fF
C685 w_n29718_2772# a_n29853_3078# 0.80fF
C686 w_n28908_3222# a_n29565_2664# 0.19fF
C687 w_n27144_n792# AlessB 0.14fF
C688 D1 adsub_b2 0.16fF
C689 a0 b0 0.82fF
C690 b3 b1 0.95fF
C691 w_n33930_n1836# a_n33840_n1809# 0.42fF
C692 w_n29898_n12546# comp_b0 2.98fF
C693 w_n29547_n10647# vdd 2.02fF
C694 comp_a2 comp_b1 0.85fF
C695 comp_b2 comp_a1 0.70fF
C696 gnd carry1 1.21fF
C697 w_n28908_5157# a_n29286_5148# 2.17fF
C698 w_n29898_n1107# a_n30123_n738# 1.20fF
C699 x3 x2 0.27fF
C700 w_n34488_n1134# vdd 2.54fF
C701 w_n33930_n1836# D 0.93fF
C702 D1 a3 0.07fF
C703 vdd x3 4.30fF
C704 a_n29880_5400# adsub_a1 1.05fF
C705 w_n29898_n1107# comp_a2 3.54fF
C706 gnd D3 4.88fF
C707 w_n31941_n14796# and_a1 0.93fF
C708 a_n30483_7947# a_n29880_7515# 1.60fF
C709 gnd a_n28998_9612# 0.60fF
C710 s0_not s0 0.07fF
C711 w_n28260_n9846# vdd 11.96fF
C712 gnd a_n30330_n2187# 0.60fF
C713 w_n29547_n1521# a_n30123_n1755# 0.66fF
C714 w_n29898_n2124# a_n30123_n1953# 0.72fF
C715 D1 adsub_b3 0.16fF
C716 w_n29547_441# vdd 2.02fF
C717 gnd comp_a0 3.10fF
C718 vdd adsub_b1 1.22fF
C719 gnd a_n30483_5832# 0.74fF
C720 w_n30402_3123# adsub_a0 0.93fF
C721 comp_a3 comp_a1 1.18fF
C722 a_n30330_n1170# a_n30123_n738# 0.99fF
C723 vdd a_n33822_n10638# 0.60fF
C724 w_n28800_n4311# a_n28710_n4284# 0.42fF
C725 w_n33462_n3807# adsub_b0 0.19fF
C726 a_n30330_n1170# comp_a2 1.80fF
C727 D a2 0.04fF
C728 carry1 sum2 0.99fF
C729 w_n35442_n12024# D1 0.19fF
C730 w_n29214_n1521# comp_a1 0.66fF
C731 w_n29898_n9288# vdd 0.48fF
C732 gnd a_n30690_7515# 0.60fF
C733 a3 b3 0.82fF
C734 w_n29898_n4491# comp_a3 1.86fF
C735 w_n33930_n396# D 0.93fF
C736 w_n29448_3528# vdd 0.48fF
C737 w_n30258_7578# adsub_b2 1.86fF
C738 w_n35442_n12024# a_n35820_n12033# 2.17fF
C739 x3 a_n28224_n6030# 0.06fF
C740 w_n30258_3528# a_n30483_3897# 1.20fF
C741 w_n28890_n7083# x3 0.84fF
C742 D1 a2 0.07fF
C743 vdd a_n33822_n8721# 0.60fF
C744 vdd a_n35820_n12888# 0.60fF
C745 gnd a_n29286_5148# 0.60fF
C746 w_n29547_n7146# vdd 1.95fF
C747 adsub_b3 w_n30258_9675# 1.86fF
C748 w_n33444_n9657# a_n33822_n9666# 2.17fF
C749 D1 adsub_a2 0.16fF
C750 vdd a_n30123_n7380# 1.04fF
C751 vdd a_n30312_9297# 0.60fF
C752 comp_b3 comp_b0 1.38fF
C753 a0 a_n33822_n9666# 0.60fF
C754 gnd AmoreB_0 1.07fF
C755 w_n35910_n12060# s1_not 0.93fF
C756 w_n29448_5463# vdd 0.48fF
C757 and_a0 and_b3 0.54fF
C758 gnd b0 3.09fF
C759 a_n30483_10044# a_n29880_9612# 1.60fF
C760 w_n30402_7173# a_n30483_7947# 0.93fF
C761 w_n29547_n10647# a_n29457_n10845# 0.19fF
C762 x2 a_n28773_n2844# 1.72fF
C763 w_n31473_n13887# and_oper_out3 0.19fF
C764 a_n29880_7515# a_n29673_7947# 0.99fF
C765 w_n28872_n5121# vdd 0.28fF
C766 x3 comp_a1 0.04fF
C767 w_n30258_5463# a_n30690_5400# 1.29fF
C768 w_n29376_3186# D1 0.93fF
C769 vdd w_n29718_8919# 2.78fF
C770 a_n30483_3897# a_n29673_3897# 0.99fF
C771 comp_a0 a_n30123_n3051# 1.27fF
C772 w_n33912_n14904# vdd 0.28fF
C773 a2 b3 0.82fF
C774 a_n33840_n1278# a1 0.60fF
C775 D1 adsub_a3 0.09fF
C776 w_n26433_n9810# a_n26811_n9819# 2.17fF
C777 w_n28260_n9846# a_n29457_n10845# 0.63fF
C778 w_n29448_7578# adsub_a2 1.86fF
C779 w_n29268_n2817# a0_not 0.19fF
C780 a_n31851_n14373# and_b2 0.60fF
C781 gnd a_n29673_5832# 1.02fF
C782 vdd adsub_a1 1.81fF
C783 w_n29178_n4194# vdd 1.86fF
C784 gnd s0 1.81fF
C785 comp_b2 a_n30123_n936# 1.98fF
C786 w_n28908_7272# a_n29565_6714# 0.19fF
C787 w_n29718_6822# a_n29853_7128# 0.80fF
C788 w_n33930_n1305# a1 0.93fF
C789 comp_a1 a_n30330_n11313# 0.60fF
C790 w_n33462_n360# a_n33840_n369# 2.17fF
C791 gnd and_a0 0.95fF
C792 w_n33912_n11079# D2 0.93fF
C793 w_n31941_n14796# and_b1 0.93fF
C794 comp_a2 a_n30123_n5067# 0.99fF
C795 w_n29898_n7749# a_n30285_n7686# 1.86fF
C796 vdd a_n29457_n8883# 1.60fF
C797 a_n30330_n7812# a_n30123_n7380# 0.99fF
C798 comp_a2 a_n30123_n9864# 0.99fF
C799 gnd a_n29880_7515# 0.60fF
C800 vdd a_n33840_n2376# 0.60fF
C801 adsub_b1 a_n30483_5634# 1.98fF
C802 w_n31473_n13887# vdd 1.14fF
C803 comp_b3 comp_b2 1.59fF
C804 w_n33912_n10170# b3 0.93fF
C805 w_n33930_n3312# vdd 0.28fF
C806 vdd D2 1.64fF
C807 a_n30483_10044# a_n29673_9846# 1.98fF
C808 gnd comp_a2 6.23fF
C809 a_n29880_9612# w_n29448_9675# 1.29fF
C810 w_n28737_n1458# comp_b1 0.63fF
C811 w_n35910_n12915# s1 0.93fF
C812 w_n35442_n12879# vdd 1.86fF
C813 comp_b0 comp_a0 0.60fF
C814 a_n29853_9225# w_n29934_9306# 0.19fF
C815 a_n30312_9297# w_n30402_9270# 0.42fF
C816 w_n28404_n756# a_n28323_n837# 0.19fF
C817 w_n29214_n5850# b1_not 0.19fF
C818 a_n29880_9612# gnd 0.60fF
C819 w_n33930_n3843# D 0.93fF
C820 w_n29547_n1521# vdd 1.95fF
C821 a_n28998_5400# carry0 2.85fF
C822 comp_b3 a_n30330_n9351# 1.06fF
C823 w_n28566_7578# carry1 1.95fF
C824 comp_a1 a_n30123_n1953# 1.98fF
C825 a_n29673_7947# a_n28998_7515# 1.08fF
C826 comp_a3 comp_b3 1.14fF
C827 w_n35910_n12501# s0_not 0.93fF
C828 w_n35910_n12060# vdd 0.28fF
C829 vdd a_n30312_3150# 0.60fF
C830 D1 a_n30483_5832# 0.99fF
C831 w_n33444_n12933# a_n33822_n12942# 2.17fF
C832 a_n30285_n7686# a_n28377_n7326# 0.06fF
C833 w_n28890_n2754# comp_b0 0.63fF
C834 w_n28872_n792# vdd 0.28fF
C835 a1 a0 0.82fF
C836 w_n28260_n9846# k 0.19fF
C837 AmoreB_0 a_n27072_n5220# 1.06fF
C838 vdd carry0 2.13fF
C839 comp_a1 a_n30123_n6282# 1.98fF
C840 a_n33840_n2871# b2 0.60fF
C841 D1 a_n30690_7515# 1.06fF
C842 w_n29205_n5004# comp_b2 0.66fF
C843 a1 a_n33822_n9135# 0.60fF
C844 w_n33462_n1800# a_n33840_n1809# 2.17fF
C845 w_n29898_n5436# a_n30123_n5265# 0.72fF
C846 w_n29547_n4833# a_n30123_n5067# 0.66fF
C847 b3 D3 0.11fF
C848 w_n29898_n11250# vdd 0.48fF
C849 w_n28737_n1458# a_n28620_n1548# 1.57fF
C850 a_n29673_9846# w_n29448_9675# 0.72fF
C851 a_n29673_10044# w_n28566_9675# 2.98fF
C852 b1 D2 0.12fF
C853 a_n30285_n7686# a_n28773_n7173# 0.80fF
C854 gnd a_n28998_7515# 0.60fF
C855 w_n29718_2772# carry0 0.14fF
C856 w_n29934_5094# a_n29853_5013# 0.19fF
C857 vdd b2 0.27fF
C858 w_n30402_5058# a_n30312_5085# 0.42fF
C859 w_n33930_n3312# b1 0.93fF
C860 w_n33930_n891# vdd 0.28fF
C861 comp_b2 comp_a0 0.39fF
C862 comp_b1 x1 0.86fF
C863 comp_b3 x3 0.62fF
C864 vdd a_n30483_3897# 0.60fF
C865 adsub_b2 adsub_a1 0.67fF
C866 w_n29547_n9630# vdd 2.02fF
C867 w_n29898_n2124# a_n30123_n1755# 1.20fF
C868 gnd a_n29457_n9828# 1.60fF
C869 D1 b0 0.19fF
C870 a_n30690_9612# adsub_b3 1.00fF
C871 w_n29898_n162# vdd 0.48fF
C872 a0 a_n33822_n13887# 0.60fF
C873 w_n29898_n3420# comp_a0 2.98fF
C874 gnd a_n30330_n3483# 0.60fF
C875 w_n29547_n11943# a_n29457_n12141# 0.19fF
C876 w_n29178_n4194# b3_not 0.19fF
C877 a2 a_n33822_n8721# 0.60fF
C878 w_n28332_n4275# a_n28710_n4284# 2.17fF
C879 vdd and_a2 0.62fF
C880 a_n28998_7515# sum2 0.99fF
C881 w_n33912_n9162# vdd 0.28fF
C882 comp_a3 comp_a0 0.49fF
C883 w_n29448_5463# a_n29673_5634# 0.72fF
C884 w_n33444_n12438# a_n33822_n12447# 2.17fF
C885 w_n28566_5463# a_n29673_5832# 2.98fF
C886 w_n33912_n15849# a_n33822_n15822# 0.42fF
C887 w_n30258_7578# a_n30690_7515# 1.29fF
C888 w_n29898_n6453# comp_b1 2.98fF
C889 w_n30258_3528# vdd 0.48fF
C890 w_n33912_n9693# a0 0.93fF
C891 adsub_b3 adsub_a1 0.67fF
C892 vdd a_n30312_7200# 0.60fF
C893 a_n29673_3897# a_n28791_3699# 1.98fF
C894 w_n29898_n9288# comp_b3 2.98fF
C895 a3 D2 0.10fF
C896 comp_a2 comp_b0 1.02fF
C897 w_n33912_n14409# a_n33822_n14382# 0.42fF
C898 w_n31473_n14364# a_n31851_n14373# 2.17fF
C899 gnd AlessB_0 1.07fF
C900 w_n29898_n7749# vdd 0.48fF
C901 vdd a_n30285_n7686# 0.02fF
C902 b2 b1 0.95fF
C903 b3 b0 0.95fF
C904 gnd a1 3.27fF
C905 a_n29673_10044# sum3 1.55fF
C906 gnd and_b2 0.60fF
C907 w_n31473_n15228# and_oper_out0 0.19fF
C908 w_n30258_5463# vdd 0.48fF
C909 sum3 w_n28566_9675# 1.20fF
C910 comp_a3 a_n28710_n4284# 0.60fF
C911 vdd a_n30123_n1755# 1.04fF
C912 w_n29898_n11250# comp_a1 1.86fF
C913 w_n33912_n15849# vdd 0.28fF
C914 adsub_a1 a_n29673_5634# 3.02fF
C915 w_n33912_n8748# a_n33822_n8721# 0.42fF
C916 a_n30483_7947# a_n29673_7749# 1.98fF
C917 w_n27576_n5085# vdd 7.49fF
C918 adsub_a3 a_n30312_9297# 1.81fF
C919 vdd a_n29673_3897# 1.21fF
C920 vdd w_n29376_9333# 0.28fF
C921 x3 comp_a0 0.41fF
C922 a_n30330_n3483# a_n30123_n3051# 0.99fF
C923 w_n27576_n5085# AmoreB 0.14fF
C924 w_n33444_n14868# vdd 1.86fF
C925 vdd a_n30123_n6084# 1.04fF
C926 w_n29448_7578# a_n29880_7515# 1.29fF
C927 w_n27144_n792# AlessB_0 1.41fF
C928 w_n29547_n3888# vdd 2.02fF
C929 vdd s1_not 0.27fF
C930 a2 D2 0.12fF
C931 comp_b2 a_n30123_n738# 0.99fF
C932 w_n33930_n1305# a_n33840_n1278# 0.42fF
C933 comp_a2 comp_b2 1.13fF
C934 w_n31941_n14796# a_n31851_n14769# 0.42fF
C935 comp_a2 a_n30330_n5499# 0.80fF
C936 w_n28890_n7083# a_n30285_n7686# 0.63fF
C937 w_n29898_n7749# a_n30330_n7812# 1.29fF
C938 a_n30330_n7812# a_n30285_n7686# 1.00fF
C939 w_n33930_n2898# b2 0.93fF
C940 w_n28566_5463# sum1 1.20fF
C941 w_n28890_n2754# x3 0.84fF
C942 w_n29178_n4194# comp_b3 0.66fF
C943 a3 b2 0.82fF
C944 adsub_b1 a_n30483_5832# 1.16fF
C945 w_n33912_n13914# vdd 0.28fF
C946 w_n35910_n12915# s0 0.93fF
C947 a_n29565_8811# w_n29718_8919# 3.02fF
C948 vdd a_n33822_n8226# 0.60fF
C949 w_n33462_n3276# vdd 1.86fF
C950 a_n30330_n12609# a_n30123_n12177# 0.99fF
C951 a_n30483_10044# a_n29673_10044# 0.99fF
C952 a_n29673_5832# a_n28791_5634# 1.98fF
C953 w_n33912_n10170# D2 0.93fF
C954 vdd a_n29565_4599# 0.60fF
C955 x2 a_n28773_n7173# 1.72fF
C956 carry2 a_n28791_9846# 1.98fF
C957 comp_a3 comp_a2 1.99fF
C958 w_n29547_n11943# vdd 2.07fF
C959 comp_a1 a_n30285_n7686# 0.04fF
C960 comp_b0 a_n30330_n3483# 1.00fF
C961 a_n30312_9297# w_n29934_9306# 2.17fF
C962 gnd x1 0.62fF
C963 w_n29898_n2124# vdd 0.48fF
C964 w_n28566_7578# a_n28998_7515# 1.29fF
C965 comp_a1 a_n30123_n1755# 1.27fF
C966 w_n33912_n8748# D2 0.93fF
C967 w_n29718_2772# a_n29637_2673# 0.96fF
C968 a_n30330_n225# comp_b3 0.60fF
C969 w_n35442_n12465# a_n35820_n12474# 2.17fF
C970 gnd a_n29286_9360# 0.60fF
C971 w_n30258_5463# a_n30483_5634# 0.72fF
C972 w_n29448_5463# a_n30483_5832# 2.98fF
C973 w_n28872_n5121# b2_not 0.93fF
C974 w_n33444_n15813# and_b0 0.19fF
C975 w_n36243_n12096# vdd 0.89fF
C976 w_n28332_54# AlessB_3 0.19fF
C977 carry2 w_n29376_9333# 0.93fF
C978 w_n33912_n14904# D3 0.93fF
C979 w_n29718_4707# a_n29565_4599# 3.02fF
C980 a2 b2 0.82fF
C981 vdd a_n33822_n15822# 0.60fF
C982 w_n27576_n756# vdd 1.86fF
C983 w_n28260_n9846# a_n28152_n9828# 1.57fF
C984 w_n33930_n891# a2 0.93fF
C985 w_n28908_3222# a_n29286_3213# 2.17fF
C986 comp_a1 a_n30123_n6084# 0.99fF
C987 gnd D0 0.60fF
C988 D a1 0.07fF
C989 a_n31851_n15237# and_b0 0.60fF
C990 w_n29898_n5436# a_n30123_n5067# 1.20fF
C991 comp_b1 a_n30123_n11079# 0.99fF
C992 w_n35910_n11592# s0_not 0.93fF
C993 a_n30330_n6516# a_n30123_n6084# 0.99fF
C994 w_n33912_n11079# vdd 0.28fF
C995 w_n28890_n7083# a_n28773_n7173# 1.57fF
C996 a_n29673_10044# w_n29448_9675# 1.20fF
C997 w_n29934_5094# a_n30312_5085# 2.17fF
C998 w_n33930_n3312# a_n33840_n3285# 0.42fF
C999 vdd a_n33840_n2871# 0.60fF
C1000 a_n30483_5832# adsub_a1 1.55fF
C1001 w_n33462_n855# vdd 1.86fF
C1002 x3 comp_a2 0.41fF
C1003 w_n29898_n1107# a_n30330_n1170# 1.29fF
C1004 gnd a_n30330_n12609# 0.60fF
C1005 w_n28890_n2754# a_n28773_n2844# 1.57fF
C1006 vdd x2 2.76fF
C1007 gnd a_n29673_10044# 1.02fF
C1008 w_n33912_n14409# b3 0.93fF
C1009 w_n33444_n11574# comp_b0 0.19fF
C1010 comp_b1 a_n28620_n1548# 0.80fF
C1011 w_n33912_n10665# a_n33822_n10638# 0.42fF
C1012 w_n29898_n10233# vdd 0.48fF
C1013 w_n28737_n1458# a1_not 0.63fF
C1014 w_n29376_5121# carry0 0.93fF
C1015 w_n35442_n12879# D3 0.19fF
C1016 w_n29718_2772# vdd 2.78fF
C1017 w_n29898_n3420# a_n30330_n3483# 1.29fF
C1018 vdd a_n33822_n10143# 0.60fF
C1019 s0 a_n35820_n12888# 0.60fF
C1020 gnd adsub_b0 1.41fF
C1021 w_n29898_n162# comp_b3 1.86fF
C1022 comp_a3 a_n30123_9# 1.98fF
C1023 adsub_a2 a_n30312_7200# 1.81fF
C1024 w_n33444_n9126# vdd 1.86fF
C1025 w_n29898_n2124# comp_a1 2.98fF
C1026 w_n29448_5463# a_n29673_5832# 1.20fF
C1027 a_n30690_3465# adsub_b0 1.00fF
C1028 w_n33444_n15813# a_n33822_n15822# 2.17fF
C1029 carry1 carry0 0.60fF
C1030 w_n29718_4707# vdd 2.78fF
C1031 w_n35442_n11556# D0 0.19fF
C1032 a1 b3 0.82fF
C1033 a3 a_n33822_n8226# 0.60fF
C1034 w_n26901_n9846# equals_d 0.93fF
C1035 temp a_n28152_n9828# 0.80fF
C1036 w_n33912_n11079# b1 0.93fF
C1037 w_n28890_n7083# x2 0.77fF
C1038 gnd a_n29853_5013# 0.60fF
C1039 w_n28890_n7083# vdd 11.51fF
C1040 D1 a_n30483_7749# 1.98fF
C1041 w_n30402_5058# adsub_b1 0.05fF
C1042 gnd a_n29286_3213# 0.60fF
C1043 comp_b0 x1 0.41fF
C1044 w_n29718_6822# vdd 2.78fF
C1045 b2 D3 0.10fF
C1046 comp_a3 a_n30123_n4320# 1.98fF
C1047 a_n29565_8811# a_n29637_8820# 1.62fF
C1048 b0 D2 0.12fF
C1049 vdd b1 0.27fF
C1050 comp_b3 a_n30285_n7686# 0.27fF
C1051 w_n33444_n15813# vdd 1.86fF
C1052 comp_b0 a_n30123_n12375# 0.99fF
C1053 adsub_a1 a_n29673_5832# 2.03fF
C1054 a_n30483_7947# a_n29673_7947# 0.99fF
C1055 w_n33444_n8712# a_n33822_n8721# 2.17fF
C1056 a_n30330_n4554# a_n30123_n4122# 0.99fF
C1057 w_n28404_n5085# vdd 1.75fF
C1058 vdd carry2 1.76fF
C1059 w_n28872_n5121# comp_a2 0.93fF
C1060 w_n29718_6822# a_n29637_6723# 0.96fF
C1061 w_n33912_n11610# D2 0.93fF
C1062 x2 comp_a1 0.04fF
C1063 w_n33444_n10629# comp_b2 0.19fF
C1064 vdd comp_a1 1.52fF
C1065 vdd w_n30402_9270# 0.28fF
C1066 vdd a_n29457_n10845# 0.80fF
C1067 gnd comp_b1 5.21fF
C1068 D1 a_n30483_9846# 1.98fF
C1069 w_n28260_n9846# a_n29457_n9828# 0.63fF
C1070 vdd a_n31851_n15237# 0.41fF
C1071 w_n31473_n14760# vdd 1.14fF
C1072 w_n29376_3186# a_n29673_3897# 0.93fF
C1073 w_n29898_n4491# vdd 0.48fF
C1074 carry0 a_n29286_5148# 1.81fF
C1075 w_n28908_7272# a_n29286_7263# 2.17fF
C1076 vdd and_a1 1.04fF
C1077 w_n33912_n10665# D2 0.93fF
C1078 gnd adsub_a0 2.13fF
C1079 w_n33930_n2898# a_n33840_n2871# 0.42fF
C1080 vdd adsub_b2 1.22fF
C1081 gnd a_n30483_7947# 0.74fF
C1082 a_n30690_5400# a_n30483_5832# 0.99fF
C1083 w_n33444_n9126# comp_a1 0.19fF
C1084 w_n27144_n792# AlessB_3 2.24fF
C1085 w_n30258_7578# a_n30483_7749# 0.72fF
C1086 w_n33444_n13878# vdd 1.86fF
C1087 comp_b0 a_n30330_n12609# 1.06fF
C1088 w_n31941_n14400# and_a2 0.93fF
C1089 comp_b2 x1 0.41fF
C1090 w_n27144_n792# AlessB_2 0.80fF
C1091 w_n28737_n5787# a_n28620_n5877# 1.57fF
C1092 gnd s0_not 0.46fF
C1093 w_n33930_n2898# vdd 0.28fF
C1094 D1 D0 0.99fF
C1095 gnd a_n30330_n1170# 0.60fF
C1096 vdd a3 0.54fF
C1097 w_n33462_n1269# a_n33840_n1278# 2.17fF
C1098 a_n30483_10044# w_n29448_9675# 2.98fF
C1099 a_n30483_9846# w_n30258_9675# 0.72fF
C1100 b2 b0 0.95fF
C1101 w_n30402_5058# adsub_a1 0.93fF
C1102 gnd a0 3.27fF
C1103 w_n28737_n1458# x3 0.81fF
C1104 w_n29718_6822# carry2 0.14fF
C1105 w_n35910_n12060# s0 1.12fF
C1106 w_n29898_n12546# vdd 0.48fF
C1107 w_n33912_n15849# D3 0.93fF
C1108 gnd a_n29286_7263# 0.60fF
C1109 a_n30483_10044# gnd 0.74fF
C1110 w_n33930_n1836# vdd 0.28fF
C1111 adsub_b3 vdd 1.22fF
C1112 a_n29673_5832# carry0 0.09fF
C1113 a_n30330_n2187# a_n30123_n1755# 0.99fF
C1114 comp_a3 x1 0.04fF
C1115 w_n30258_5463# a_n30483_5832# 1.20fF
C1116 w_n28872_n5121# a_n28782_n5094# 0.42fF
C1117 w_n31941_n15264# and_b0 0.93fF
C1118 w_n35442_n12024# vdd 1.86fF
C1119 AlessB_0 a_n27072_n891# 1.06fF
C1120 w_n33930_n2403# D 0.93fF
C1121 w_n28404_n756# vdd 1.75fF
C1122 w_n29448_7578# a_n29673_7749# 0.72fF
C1123 w_n33912_n10665# b2 0.93fF
C1124 w_n29934_3159# a_n29853_3078# 0.19fF
C1125 w_n30402_3123# a_n30312_3150# 0.42fF
C1126 w_n33444_n14373# and_b3 0.19fF
C1127 D1 adsub_b0 0.45fF
C1128 comp_a1 a_n30330_n6516# 1.77fF
C1129 comp_b2 a_n28782_n765# 0.60fF
C1130 w_n33462_n855# adsub_a2 0.19fF
C1131 w_n29898_n5436# comp_b2 3.54fF
C1132 w_n29898_n5436# a_n30330_n5499# 1.29fF
C1133 vdd a2 1.14fF
C1134 comp_b1 a_n30123_n10881# 1.27fF
C1135 w_n35910_n11592# a_n35820_n11565# 0.42fF
C1136 gnd and_b3 0.60fF
C1137 w_n33444_n11043# vdd 1.86fF
C1138 comp_b2 a_n30123_n5265# 1.98fF
C1139 w_n33912_n13914# D3 0.93fF
C1140 gnd a_n29673_7947# 1.02fF
C1141 vdd adsub_a2 1.81fF
C1142 w_n33462_n3276# a_n33840_n3285# 2.17fF
C1143 a_n29880_3465# adsub_a0 1.05fF
C1144 comp_b2 a_n30123_n10062# 0.99fF
C1145 a3 b1 0.82fF
C1146 w_n33930_n1305# D 0.93fF
C1147 a_n30483_5832# a_n29880_5400# 1.60fF
C1148 w_n33930_n396# vdd 0.28fF
C1149 D1 a_n29286_3213# 1.81fF
C1150 w_n33444_n10629# a_n33822_n10638# 2.17fF
C1151 w_n33912_n10170# vdd 0.28fF
C1152 comp_b0 comp_b1 0.98fF
C1153 x3 x1 0.27fF
C1154 w_n33912_n15849# b0 0.93fF
C1155 comp_b3 x2 0.41fF
C1156 w_n27576_n5085# AmoreB_0 1.41fF
C1157 vdd and_b1 1.06fF
C1158 vdd comp_b3 2.00fF
C1159 w_n29376_3186# vdd 0.28fF
C1160 comp_b0 a_n30123_n3249# 1.98fF
C1161 w_n30402_3123# a_n30483_3897# 0.93fF
C1162 adsub_a3 vdd 1.81fF
C1163 carry0 sum1 0.99fF
C1164 gnd a_n30690_3465# 0.60fF
C1165 w_n33912_n10170# a_n33822_n10143# 0.42fF
C1166 a_n29673_7947# sum2 1.55fF
C1167 comp_a3 a_n30123_207# 1.27fF
C1168 w_n33912_n8748# vdd 0.28fF
C1169 w_n29898_n2124# a_n30330_n2187# 1.29fF
C1170 adsub_b3 w_n30402_9270# 0.05fF
C1171 vdd a_n29565_8811# 0.60fF
C1172 w_n33930_n2403# b3 0.93fF
C1173 w_n28044_n5121# a_n27954_n5094# 0.42fF
C1174 w_n29376_5121# vdd 0.28fF
C1175 AmoreB_3 a_n27072_n5220# 1.04fF
C1176 w_n28872_n792# a2_not 0.93fF
C1177 comp_a3 a_n30123_n9117# 1.98fF
C1178 a_n33840_n1809# a0 0.60fF
C1179 a2 b1 0.82fF
C1180 w_n34488_n1134# D0 0.80fF
C1181 a_n29457_n12141# a_n28152_n9828# 0.80fF
C1182 gnd a_n30330_n4554# 0.60fF
C1183 w_n33444_n14373# a_n33822_n14382# 2.17fF
C1184 D1 adsub_a0 0.07fF
C1185 w_n29214_n5850# vdd 1.29fF
C1186 vdd a_n33822_n11583# 0.60fF
C1187 D1 a_n30483_7947# 0.99fF
C1188 a1 D2 0.12fF
C1189 comp_a2 a_n30285_n7686# 0.27fF
C1190 D a0 0.07fF
C1191 w_n29376_7236# vdd 0.28fF
C1192 comp_a3 a_n30123_n4122# 0.99fF
C1193 comp_b2 comp_b1 2.24fF
C1194 vdd carry1 1.27fF
C1195 vdd a_n33840_n3285# 0.60fF
C1196 vdd a_n28710_45# 0.41fF
C1197 a_n29880_5400# a_n29673_5832# 0.99fF
C1198 w_n31941_n15264# vdd 0.28fF
C1199 w_n29898_n1107# comp_b2 1.86fF
C1200 comp_b0 a_n30123_n12177# 1.27fF
C1201 gnd and_a3 0.66fF
C1202 a_n29565_2664# a_n29637_2673# 1.62fF
C1203 s1_not s0 0.04fF
C1204 w_n29205_n5004# vdd 1.92fF
C1205 w_n29268_n7146# b0_not 0.19fF
C1206 vdd w_n29934_9306# 1.86fF
C1207 vdd a_n26811_n9819# 0.41fF
C1208 x3 a_n28224_n1701# 0.06fF
C1209 x1 a_n28773_n2844# 1.58fF
C1210 D1 a_n30483_10044# 0.99fF
C1211 vdd a_n33822_n15291# 0.60fF
C1212 w_n31941_n14400# vdd 0.28fF
C1213 w_n29547_n9630# a_n29457_n9828# 0.19fF
C1214 w_n29448_7578# a_n30483_7947# 2.98fF
C1215 x2 comp_a0 0.41fF
C1216 w_n29898_n3420# a_n30123_n3249# 0.72fF
C1217 w_n29547_n2817# a_n30123_n3051# 0.66fF
C1218 vdd comp_a0 0.96fF
C1219 w_n28566_3528# sum0 1.20fF
C1220 vdd a_n30483_5832# 0.60fF
C1221 comp_b3 comp_a1 1.61fF
C1222 w_n33930_n3843# vdd 0.28fF
C1223 comp_a3 comp_b1 0.65fF
C1224 w_n29718_4707# carry1 0.14fF
C1225 a_n30330_n1170# comp_b2 0.60fF
C1226 w_n30402_7173# a_n30312_7200# 0.42fF
C1227 a3 a2 0.82fF
C1228 w_n29934_7209# a_n29853_7128# 0.19fF
C1229 w_n28332_n4275# AmoreB_3 0.19fF
C1230 vdd a_n33822_n13356# 0.60fF
C1231 w_n33912_n14904# a_n33822_n14877# 0.42fF
C1232 gnd a_n29880_3465# 0.60fF
C1233 carry1 a_n28791_7749# 1.98fF
C1234 w_n29898_n162# a_n30123_9# 0.72fF
C1235 w_n29547_441# a_n30123_207# 0.66fF
C1236 adsub_a3 w_n30402_9270# 0.93fF
C1237 w_n33444_n12438# and_a3 0.19fF
C1238 adsub_b0 a_n30483_3699# 1.98fF
C1239 b0 a_n33822_n15822# 0.60fF
C1240 w_n29898_n4491# comp_b3 2.98fF
C1241 w_n33912_n13383# vdd 0.28fF
C1242 w_n33930_n396# a3 0.93fF
C1243 w_n30258_7578# a_n30483_7947# 1.20fF
C1244 and_a1 and_b1 2.13fF
C1245 w_n28890_n2754# x2 0.77fF
C1246 a_n33822_n15822# Gnd 6.54fF
C1247 and_oper_out0 Gnd 0.88fF
C1248 and_b0 Gnd 33.08fF
C1249 a_n31851_n15237# Gnd 6.54fF
C1250 a_n33822_n15291# Gnd 6.54fF
C1251 and_oper_out1 Gnd 0.88fF
C1252 and_b1 Gnd 31.42fF
C1253 a_n31851_n14769# Gnd 6.54fF
C1254 a_n33822_n14877# Gnd 6.54fF
C1255 and_oper_out2 Gnd 0.88fF
C1256 and_b2 Gnd 30.06fF
C1257 a_n31851_n14373# Gnd 6.54fF
C1258 a_n33822_n14382# Gnd 6.54fF
C1259 and_oper_out3 Gnd 0.88fF
C1260 and_b3 Gnd 30.52fF
C1261 a_n31851_n13896# Gnd 6.54fF
C1262 and_a0 Gnd 14.31fF
C1263 a_n33822_n13887# Gnd 6.54fF
C1264 and_a1 Gnd 12.22fF
C1265 a_n33822_n13356# Gnd 6.54fF
C1266 and_a2 Gnd 12.81fF
C1267 a_n33822_n12942# Gnd 6.54fF
C1268 a_n30123_n12375# Gnd 11.04fF
C1269 a_n30123_n12177# Gnd 16.56fF
C1270 a_n35820_n12888# Gnd 6.54fF
C1271 and_a3 Gnd 13.30fF
C1272 D3 Gnd 137.57fF
C1273 a_n33822_n12447# Gnd 6.54fF
C1274 a_n30330_n12609# Gnd 43.58fF
C1275 s1 Gnd 35.20fF
C1276 a_n35820_n12474# Gnd 6.54fF
C1277 a_n30123_n11079# Gnd 11.04fF
C1278 a_n30123_n10881# Gnd 16.56fF
C1279 a_n30330_n11313# Gnd 43.58fF
C1280 AequalsB Gnd 0.88fF
C1281 equals_d Gnd 1.86fF
C1282 k Gnd 16.19fF
C1283 a_n28152_n9828# Gnd 11.33fF
C1284 temp Gnd 2.34fF
C1285 a_n29457_n12141# Gnd 86.30fF
C1286 a_n29457_n10845# Gnd 58.33fF
C1287 a_n26811_n9819# Gnd 6.54fF
C1288 a_n29457_n9828# Gnd 48.53fF
C1289 a_n30123_n10062# Gnd 11.04fF
C1290 a_n30123_n9864# Gnd 16.56fF
C1291 a_n30330_n10296# Gnd 43.58fF
C1292 a_n29457_n8883# Gnd 64.10fF
C1293 a_n30123_n9117# Gnd 11.04fF
C1294 a_n30123_n8919# Gnd 16.56fF
C1295 a_n30330_n9351# Gnd 43.58fF
C1296 a_n29457_n7344# Gnd 0.88fF
C1297 a_n28773_n7173# Gnd 11.33fF
C1298 b0_not Gnd 7.18fF
C1299 a_n30123_n7578# Gnd 10.80fF
C1300 a_n30123_n7380# Gnd 16.56fF
C1301 a_n30285_n7686# Gnd 36.63fF
C1302 a_n30330_n7812# Gnd 43.58fF
C1303 a_n33822_n11583# Gnd 6.54fF
C1304 a_n33822_n11052# Gnd 6.54fF
C1305 a_n35820_n12033# Gnd 6.54fF
C1306 s0 Gnd 61.18fF
C1307 s1_not Gnd 11.65fF
C1308 s0_not Gnd 21.63fF
C1309 a_n35820_n11565# Gnd 6.54fF
C1310 a_n33822_n10638# Gnd 6.54fF
C1311 a_n33822_n10143# Gnd 6.54fF
C1312 a_n33822_n9666# Gnd 6.54fF
C1313 a_n33822_n9135# Gnd 6.54fF
C1314 a_n33822_n8721# Gnd 6.54fF
C1315 a_n28620_n5877# Gnd 11.33fF
C1316 temp_more Gnd 2.93fF
C1317 b1_not Gnd 8.22fF
C1318 a_n30123_n6282# Gnd 10.80fF
C1319 a_n30123_n6084# Gnd 16.56fF
C1320 a_n30330_n6516# Gnd 43.58fF
C1321 AmoreB Gnd 0.76fF
C1322 a_n27072_n5220# Gnd 5.08fF
C1323 AmoreB_0 Gnd 34.46fF
C1324 AmoreB_1 Gnd 20.13fF
C1325 AmoreB_2 Gnd 5.74fF
C1326 a_n27954_n5094# Gnd 6.40fF
C1327 a_n28323_n5166# Gnd 11.54fF
C1328 b2_not Gnd 9.42fF
C1329 a_n28782_n5094# Gnd 6.54fF
C1330 a_n30123_n5265# Gnd 10.80fF
C1331 a_n30123_n5067# Gnd 16.56fF
C1332 a_n30330_n5499# Gnd 43.58fF
C1333 AmoreB_3 Gnd 29.29fF
C1334 b3_not Gnd 10.81fF
C1335 a_n28710_n4284# Gnd 6.54fF
C1336 a_n30123_n4320# Gnd 10.80fF
C1337 a_n30123_n4122# Gnd 16.56fF
C1338 a_n30330_n4554# Gnd 43.58fF
C1339 x0 Gnd 0.88fF
C1340 a_n28773_n2844# Gnd 11.33fF
C1341 a0_not Gnd 7.18fF
C1342 a_n30123_n3249# Gnd 10.80fF
C1343 a_n30123_n3051# Gnd 16.56fF
C1344 comp_a0 Gnd 186.07fF
C1345 a_n30330_n3483# Gnd 43.58fF
C1346 x1 Gnd 36.32fF
C1347 a_n28620_n1548# Gnd 11.33fF
C1348 temp_less Gnd 2.93fF
C1349 a1_not Gnd 8.22fF
C1350 a_n30123_n1953# Gnd 10.80fF
C1351 a_n30123_n1755# Gnd 16.56fF
C1352 comp_b1 Gnd 416.68fF
C1353 comp_a1 Gnd 307.44fF
C1354 a_n30330_n2187# Gnd 43.58fF
C1355 AlessB Gnd 0.76fF
C1356 a_n27072_n891# Gnd 5.08fF
C1357 AlessB_0 Gnd 34.46fF
C1358 AlessB_1 Gnd 20.13fF
C1359 AlessB_2 Gnd 5.74fF
C1360 a_n27954_n765# Gnd 6.40fF
C1361 a_n28323_n837# Gnd 11.54fF
C1362 a2_not Gnd 9.42fF
C1363 a_n28782_n765# Gnd 6.54fF
C1364 x2 Gnd 51.94fF
C1365 a_n30123_n936# Gnd 10.80fF
C1366 a_n30123_n738# Gnd 16.56fF
C1367 D2 Gnd 152.21fF
C1368 a_n33822_n8226# Gnd 6.54fF
C1369 comp_b0 Gnd 337.58fF
C1370 b0 Gnd 87.79fF
C1371 a_n33840_n3816# Gnd 6.54fF
C1372 b1 Gnd 83.59fF
C1373 a_n33840_n3285# Gnd 6.54fF
C1374 b2 Gnd 75.06fF
C1375 a_n33840_n2871# Gnd 6.54fF
C1376 b3 Gnd 71.29fF
C1377 a_n33840_n2376# Gnd 6.54fF
C1378 a0 Gnd 91.84fF
C1379 a_n33840_n1809# Gnd 6.54fF
C1380 a1 Gnd 91.61fF
C1381 a_n33840_n1278# Gnd 6.54fF
C1382 a_n34407_n1233# Gnd 3.59fF
C1383 D0 Gnd 313.55fF
C1384 a_n33840_n864# Gnd 6.54fF
C1385 a2 Gnd 73.93fF
C1386 comp_b2 Gnd 327.30fF
C1387 comp_a2 Gnd 294.37fF
C1388 a_n30330_n1170# Gnd 43.58fF
C1389 a3 Gnd 71.74fF
C1390 D Gnd 106.69fF
C1391 AlessB_3 Gnd 29.29fF
C1392 a3_not Gnd 10.81fF
C1393 a_n28710_45# Gnd 6.54fF
C1394 x3 Gnd 73.38fF
C1395 a_n30123_9# Gnd 10.80fF
C1396 a_n30123_207# Gnd 16.56fF
C1397 a_n33840_n369# Gnd 6.54fF
C1398 comp_b3 Gnd 315.86fF
C1399 comp_a3 Gnd 375.69fF
C1400 a_n30330_n225# Gnd 43.58fF
C1401 a_n29637_2673# Gnd 3.38fF
C1402 a_n29565_2664# Gnd 26.35fF
C1403 a_n29286_3213# Gnd 6.13fF
C1404 a_n29853_3078# Gnd 13.17fF
C1405 a_n30312_3150# Gnd 6.26fF
C1406 a_n28791_3699# Gnd 10.80fF
C1407 sum0 Gnd 12.42fF
C1408 a_n28998_3465# Gnd 43.33fF
C1409 a_n29673_3699# Gnd 10.80fF
C1410 a_n29673_3897# Gnd 63.56fF
C1411 adsub_a0 Gnd 185.44fF
C1412 a_n29880_3465# Gnd 43.33fF
C1413 a_n30483_3699# Gnd 10.80fF
C1414 a_n30483_3897# Gnd 66.86fF
C1415 adsub_b0 Gnd 71.70fF
C1416 a_n30690_3465# Gnd 43.58fF
C1417 a_n29637_4608# Gnd 3.38fF
C1418 a_n29565_4599# Gnd 26.35fF
C1419 a_n29286_5148# Gnd 6.13fF
C1420 a_n29853_5013# Gnd 13.17fF
C1421 a_n30312_5085# Gnd 6.26fF
C1422 a_n28791_5634# Gnd 10.80fF
C1423 sum1 Gnd 12.42fF
C1424 carry0 Gnd 85.53fF
C1425 a_n28998_5400# Gnd 43.33fF
C1426 a_n29673_5634# Gnd 10.80fF
C1427 a_n29673_5832# Gnd 63.56fF
C1428 adsub_a1 Gnd 211.31fF
C1429 a_n29880_5400# Gnd 43.33fF
C1430 a_n30483_5634# Gnd 10.80fF
C1431 a_n30483_5832# Gnd 66.86fF
C1432 adsub_b1 Gnd 54.50fF
C1433 a_n30690_5400# Gnd 43.58fF
C1434 a_n29637_6723# Gnd 3.38fF
C1435 a_n29565_6714# Gnd 26.35fF
C1436 a_n29286_7263# Gnd 6.13fF
C1437 a_n29853_7128# Gnd 13.17fF
C1438 a_n30312_7200# Gnd 6.26fF
C1439 a_n28791_7749# Gnd 10.80fF
C1440 sum2 Gnd 12.42fF
C1441 carry1 Gnd 141.82fF
C1442 a_n28998_7515# Gnd 43.33fF
C1443 a_n29673_7749# Gnd 10.80fF
C1444 a_n29673_7947# Gnd 63.56fF
C1445 adsub_a2 Gnd 224.19fF
C1446 a_n29880_7515# Gnd 43.33fF
C1447 a_n30483_7749# Gnd 10.80fF
C1448 a_n30483_7947# Gnd 66.86fF
C1449 adsub_b2 Gnd 58.25fF
C1450 a_n30690_7515# Gnd 43.58fF
C1451 carry3 Gnd 0.76fF
C1452 a_n29637_8820# Gnd 3.38fF
C1453 a_n29565_8811# Gnd 26.35fF
C1454 a_n29286_9360# Gnd 6.13fF
C1455 a_n29853_9225# Gnd 13.17fF
C1456 a_n30312_9297# Gnd 6.26fF
C1457 a_n28791_9846# Gnd 10.80fF
C1458 sum3 Gnd 12.42fF
C1459 carry2 Gnd 131.59fF
C1460 a_n28998_9612# Gnd 43.33fF
C1461 a_n29673_9846# Gnd 10.80fF
C1462 a_n29673_10044# Gnd 63.56fF
C1463 vdd Gnd 1103.38fF
C1464 gnd Gnd 1551.22fF
C1465 adsub_a3 Gnd 245.84fF
C1466 a_n29880_9612# Gnd 43.33fF
C1467 a_n30483_9846# Gnd 10.80fF
C1468 a_n30483_10044# Gnd 66.86fF
C1469 adsub_b3 Gnd 61.87fF
C1470 D1 Gnd 980.84fF
C1471 a_n30690_9612# Gnd 43.58fF
C1472 w_n33912_n15849# Gnd 29.29fF
C1473 w_n33444_n15813# Gnd 28.07fF
C1474 w_n31941_n15264# Gnd 29.29fF
C1475 w_n33912_n15318# Gnd 29.29fF
C1476 w_n33444_n15282# Gnd 28.07fF
C1477 w_n31473_n15228# Gnd 28.07fF
C1478 w_n31941_n14796# Gnd 29.29fF
C1479 w_n33912_n14904# Gnd 29.29fF
C1480 w_n33444_n14868# Gnd 28.07fF
C1481 w_n31473_n14760# Gnd 28.07fF
C1482 w_n31941_n14400# Gnd 29.29fF
C1483 w_n33912_n14409# Gnd 29.29fF
C1484 w_n31473_n14364# Gnd 28.07fF
C1485 w_n33444_n14373# Gnd 28.07fF
C1486 w_n31941_n13923# Gnd 29.29fF
C1487 w_n31473_n13887# Gnd 28.07fF
C1488 w_n33912_n13914# Gnd 29.29fF
C1489 w_n33444_n13878# Gnd 28.07fF
C1490 w_n33912_n13383# Gnd 29.29fF
C1491 w_n33444_n13347# Gnd 28.07fF
C1492 w_n33912_n12969# Gnd 29.29fF
C1493 w_n33444_n12933# Gnd 28.07fF
C1494 w_n35910_n12915# Gnd 29.29fF
C1495 w_n35442_n12879# Gnd 28.07fF
C1496 w_n29547_n11943# Gnd 26.52fF
C1497 w_n29898_n12546# Gnd 73.22fF
C1498 w_n33912_n12474# Gnd 29.29fF
C1499 w_n35910_n12501# Gnd 29.29fF
C1500 w_n36234_n12420# Gnd 28.47fF
C1501 w_n33444_n12438# Gnd 28.07fF
C1502 w_n35442_n12465# Gnd 28.07fF
C1503 w_n35910_n12060# Gnd 29.29fF
C1504 w_n36243_n12096# Gnd 24.41fF
C1505 w_n35442_n12024# Gnd 28.07fF
C1506 w_n33912_n11610# Gnd 29.29fF
C1507 w_n33444_n11574# Gnd 28.07fF
C1508 w_n35910_n11592# Gnd 29.29fF
C1509 w_n35442_n11556# Gnd 28.07fF
C1510 w_n29547_n10647# Gnd 26.36fF
C1511 w_n29898_n11250# Gnd 73.22fF
C1512 w_n33912_n11079# Gnd 29.29fF
C1513 w_n33444_n11043# Gnd 28.07fF
C1514 w_n33912_n10665# Gnd 29.29fF
C1515 w_n33444_n10629# Gnd 28.07fF
C1516 w_n26901_n9846# Gnd 29.29fF
C1517 w_n26433_n9810# Gnd 28.07fF
C1518 w_n28260_n9846# Gnd 161.09fF
C1519 w_n29547_n9630# Gnd 26.36fF
C1520 w_n29898_n10233# Gnd 73.22fF
C1521 w_n33912_n10170# Gnd 29.29fF
C1522 w_n33444_n10134# Gnd 28.07fF
C1523 w_n33912_n9693# Gnd 29.29fF
C1524 w_n33444_n9657# Gnd 28.07fF
C1525 w_n29547_n8685# Gnd 26.36fF
C1526 w_n29898_n9288# Gnd 73.22fF
C1527 w_n33912_n9162# Gnd 29.29fF
C1528 w_n33444_n9126# Gnd 28.07fF
C1529 w_n33912_n8748# Gnd 29.29fF
C1530 w_n33444_n8712# Gnd 28.07fF
C1531 w_n33912_n8253# Gnd 29.29fF
C1532 w_n33444_n8217# Gnd 28.07fF
C1533 w_n29268_n7146# Gnd 26.36fF
C1534 w_n29547_n7146# Gnd 25.95fF
C1535 w_n29898_n7749# Gnd 73.22fF
C1536 w_n28890_n7083# Gnd 161.33fF
C1537 w_n29214_n5850# Gnd 26.36fF
C1538 w_n29547_n5850# Gnd 25.95fF
C1539 w_n29898_n6453# Gnd 73.22fF
C1540 w_n28737_n5787# Gnd 161.33fF
C1541 w_n28044_n5121# Gnd 29.29fF
C1542 w_n28872_n5121# Gnd 29.29fF
C1543 w_n27576_n5085# Gnd 95.92fF
C1544 w_n28404_n5085# Gnd 28.07fF
C1545 w_n29205_n5004# Gnd 26.52fF
C1546 w_n29547_n4833# Gnd 26.36fF
C1547 w_n29898_n5436# Gnd 73.22fF
C1548 w_n28800_n4311# Gnd 29.29fF
C1549 w_n28332_n4275# Gnd 28.07fF
C1550 w_n29178_n4194# Gnd 26.36fF
C1551 w_n29547_n3888# Gnd 26.36fF
C1552 w_n29898_n4491# Gnd 73.22fF
C1553 w_n33930_n3843# Gnd 29.29fF
C1554 w_n33462_n3807# Gnd 28.07fF
C1555 w_n29268_n2817# Gnd 26.36fF
C1556 w_n29547_n2817# Gnd 25.95fF
C1557 w_n29898_n3420# Gnd 73.22fF
C1558 w_n33930_n3312# Gnd 29.29fF
C1559 w_n33462_n3276# Gnd 28.07fF
C1560 w_n33930_n2898# Gnd 29.29fF
C1561 w_n28890_n2754# Gnd 161.33fF
C1562 w_n33462_n2862# Gnd 28.07fF
C1563 w_n33930_n2403# Gnd 29.29fF
C1564 w_n33462_n2367# Gnd 28.07fF
C1565 w_n29214_n1521# Gnd 26.36fF
C1566 w_n29547_n1521# Gnd 25.95fF
C1567 w_n29898_n2124# Gnd 73.22fF
C1568 w_n33930_n1836# Gnd 29.29fF
C1569 w_n33462_n1800# Gnd 28.07fF
C1570 w_n28737_n1458# Gnd 161.33fF
C1571 w_n33930_n1305# Gnd 29.29fF
C1572 w_n27144_n792# Gnd 62.16fF
C1573 w_n28044_n792# Gnd 29.29fF
C1574 w_n28872_n792# Gnd 29.29fF
C1575 w_n27576_n756# Gnd 28.07fF
C1576 w_n28404_n756# Gnd 28.07fF
C1577 w_n29205_n675# Gnd 26.52fF
C1578 w_n29547_n504# Gnd 26.36fF
C1579 w_n29898_n1107# Gnd 73.22fF
C1580 w_n33462_n1269# Gnd 28.07fF
C1581 w_n34488_n1134# Gnd 41.25fF
C1582 w_n33930_n891# Gnd 29.29fF
C1583 w_n33462_n855# Gnd 28.07fF
C1584 w_n33930_n396# Gnd 29.29fF
C1585 w_n33462_n360# Gnd 28.07fF
C1586 w_n28800_18# Gnd 29.29fF
C1587 w_n28332_54# Gnd 28.07fF
C1588 w_n29178_135# Gnd 26.36fF
C1589 w_n29547_441# Gnd 26.36fF
C1590 w_n29898_n162# Gnd 73.22fF
C1591 w_n29718_2772# Gnd 41.25fF
C1592 w_n29376_3186# Gnd 29.29fF
C1593 w_n30402_3123# Gnd 29.29fF
C1594 w_n29934_3159# Gnd 28.07fF
C1595 w_n28908_3222# Gnd 28.07fF
C1596 w_n28566_3528# Gnd 73.22fF
C1597 w_n29448_3528# Gnd 73.22fF
C1598 w_n30258_3528# Gnd 73.22fF
C1599 w_n29718_4707# Gnd 41.25fF
C1600 w_n29376_5121# Gnd 29.29fF
C1601 w_n30402_5058# Gnd 29.29fF
C1602 w_n29934_5094# Gnd 28.07fF
C1603 w_n28908_5157# Gnd 28.07fF
C1604 w_n28566_5463# Gnd 73.22fF
C1605 w_n29448_5463# Gnd 73.22fF
C1606 w_n30258_5463# Gnd 73.22fF
C1607 w_n29718_6822# Gnd 41.25fF
C1608 w_n29376_7236# Gnd 29.29fF
C1609 w_n30402_7173# Gnd 29.29fF
C1610 w_n29934_7209# Gnd 28.07fF
C1611 w_n28908_7272# Gnd 28.07fF
C1612 w_n28566_7578# Gnd 73.22fF
C1613 w_n29448_7578# Gnd 73.22fF
C1614 w_n30258_7578# Gnd 73.22fF
C1615 w_n29718_8919# Gnd 41.25fF
C1616 w_n29376_9333# Gnd 29.29fF
C1617 w_n30402_9270# Gnd 29.29fF
C1618 w_n29934_9306# Gnd 28.07fF
C1619 w_n28908_9369# Gnd 28.07fF
C1620 w_n28566_9675# Gnd 73.22fF
C1621 w_n29448_9675# Gnd 73.22fF
C1622 w_n30258_9675# Gnd 73.22fF




.tran 0.1n 400n

.measure tran trise 
+ TRIG v(A1) VAL = 'SUPPLY/2' TD = 0ns RISE =1 
+ TARG v(AmoreB) VAL = 'SUPPLY/2' TD = 0ns RISE =1S

.measure tran tfall 
+ TRIG v(A1) VAL = 'SUPPLY/2' TD = 0ns FALL =1 
+ TARG v(AmoreB) VAL = 'SUPPLY/2' TD = 0ns FALL=1 

.measure tran tpd param = '(trise + tfall)/2' goal = 0
        
.control
run 
plot v(s0) v(s1)+2
plot v(D0) v(D1)+2 v(D2)+4 v(D3)+6
plot v(a0) v(a1)+2 v(a2)+4 v(a3)+6
plot v(b0) v(b1)+2 v(b2)+4 v(b3)+6

plot v(and_a0) v(and_a1)+2 v(and_a2)+4 v(and_a3)+6
plot v(and_b0) v(and_b1)+2 v(and_b2)+4 v(and_b3)+6

plot v(comp_a0) v(comp_a1)+2 v(comp_a2)+4 v(comp_a3)+6
plot v(comp_b0) v(comp_b1)+2 v(comp_b2)+4 v(comp_b3)+6

plot v(adsub_a0) v(adsub_a1)+2 v(adsub_a2)+4 v(adsub_a3)+6
plot v(adsub_b0) v(adsub_b1)+2 v(adsub_b2)+4 v(adsub_b3)+6

plot v(and_oper_out3)+8 v(and_oper_out2)+6 v(and_oper_out1)+4 v(and_oper_out0)+2

plot v(AmoreB) v(AlessB)+2 v(AequalsB)+4

plot v(sum0) v(sum1)+2 v(sum2)+4 v(sum3)+6 v(carry3)+8
quit
.endc
.endc