magic
tech scmos
magscale 9 1
timestamp 1700920797
<< nwell >>
rect 220 71 241 77
rect 168 54 204 64
rect 220 59 237 71
rect 220 58 227 59
rect 229 58 237 59
rect 220 16 241 22
rect 168 -1 204 9
rect 220 4 237 16
rect 220 3 227 4
rect 229 3 237 4
rect 106 -28 145 -15
rect 220 -30 241 -24
rect 168 -47 204 -37
rect 220 -42 237 -30
rect 220 -43 227 -42
rect 229 -43 237 -42
rect 220 -89 241 -83
rect 168 -106 204 -96
rect 220 -101 237 -89
rect 220 -102 227 -101
rect 229 -102 237 -101
rect 220 -152 241 -146
rect 168 -169 204 -159
rect 220 -164 237 -152
rect 220 -165 227 -164
rect 229 -165 237 -164
rect 220 -207 241 -201
rect 168 -224 204 -214
rect 220 -219 237 -207
rect 220 -220 227 -219
rect 229 -220 237 -219
rect 220 -253 241 -247
rect 168 -270 204 -260
rect 220 -265 237 -253
rect 220 -266 227 -265
rect 229 -266 237 -265
rect 220 -312 241 -306
rect 168 -329 204 -319
rect 220 -324 237 -312
rect 220 -325 227 -324
rect 229 -325 237 -324
<< ntransistor >>
rect 227 49 229 52
rect 176 43 178 46
rect 194 43 196 46
rect 227 -6 229 -3
rect 176 -12 178 -9
rect 194 -12 196 -9
rect 113 -39 115 -36
rect 123 -39 125 -36
rect 137 -39 139 -36
rect 227 -52 229 -49
rect 176 -58 178 -55
rect 194 -58 196 -55
rect 227 -111 229 -108
rect 176 -117 178 -114
rect 194 -117 196 -114
rect 227 -174 229 -171
rect 176 -180 178 -177
rect 194 -180 196 -177
rect 227 -229 229 -226
rect 176 -235 178 -232
rect 194 -235 196 -232
rect 227 -275 229 -272
rect 176 -281 178 -278
rect 194 -281 196 -278
rect 227 -334 229 -331
rect 176 -340 178 -337
rect 194 -340 196 -337
<< ptransistor >>
rect 176 57 178 62
rect 194 57 196 62
rect 227 60 229 66
rect 176 2 178 7
rect 194 2 196 7
rect 227 5 229 11
rect 113 -26 115 -21
rect 123 -26 125 -21
rect 137 -26 139 -21
rect 176 -44 178 -39
rect 194 -44 196 -39
rect 227 -41 229 -35
rect 176 -103 178 -98
rect 194 -103 196 -98
rect 227 -100 229 -94
rect 176 -166 178 -161
rect 194 -166 196 -161
rect 227 -163 229 -157
rect 176 -221 178 -216
rect 194 -221 196 -216
rect 227 -218 229 -212
rect 176 -267 178 -262
rect 194 -267 196 -262
rect 227 -264 229 -258
rect 176 -326 178 -321
rect 194 -326 196 -321
rect 227 -323 229 -317
<< ndiffusion >>
rect 222 51 227 52
rect 222 49 223 51
rect 226 49 227 51
rect 229 49 231 52
rect 234 49 235 52
rect 172 45 176 46
rect 172 43 173 45
rect 175 43 176 45
rect 178 43 194 46
rect 196 44 197 46
rect 199 44 200 46
rect 196 43 200 44
rect 222 -4 227 -3
rect 222 -6 223 -4
rect 226 -6 227 -4
rect 229 -6 231 -3
rect 234 -6 235 -3
rect 172 -10 176 -9
rect 172 -12 173 -10
rect 175 -12 176 -10
rect 178 -12 194 -9
rect 196 -11 197 -9
rect 199 -11 200 -9
rect 196 -12 200 -11
rect 109 -38 110 -36
rect 112 -38 113 -36
rect 109 -39 113 -38
rect 115 -38 116 -36
rect 115 -39 118 -38
rect 119 -38 120 -36
rect 122 -38 123 -36
rect 119 -39 123 -38
rect 125 -38 126 -36
rect 125 -39 128 -38
rect 133 -38 134 -36
rect 136 -38 137 -36
rect 133 -39 137 -38
rect 139 -38 140 -36
rect 142 -38 143 -36
rect 139 -39 143 -38
rect 222 -50 227 -49
rect 222 -52 223 -50
rect 226 -52 227 -50
rect 229 -52 231 -49
rect 234 -52 235 -49
rect 172 -56 176 -55
rect 172 -58 173 -56
rect 175 -58 176 -56
rect 178 -58 194 -55
rect 196 -57 197 -55
rect 199 -57 200 -55
rect 196 -58 200 -57
rect 222 -109 227 -108
rect 222 -111 223 -109
rect 226 -111 227 -109
rect 229 -111 231 -108
rect 234 -111 235 -108
rect 172 -115 176 -114
rect 172 -117 173 -115
rect 175 -117 176 -115
rect 178 -117 194 -114
rect 196 -116 197 -114
rect 199 -116 200 -114
rect 196 -117 200 -116
rect 222 -172 227 -171
rect 222 -174 223 -172
rect 226 -174 227 -172
rect 229 -174 231 -171
rect 234 -174 235 -171
rect 172 -178 176 -177
rect 172 -180 173 -178
rect 175 -180 176 -178
rect 178 -180 194 -177
rect 196 -179 197 -177
rect 199 -179 200 -177
rect 196 -180 200 -179
rect 222 -227 227 -226
rect 222 -229 223 -227
rect 226 -229 227 -227
rect 229 -229 231 -226
rect 234 -229 235 -226
rect 172 -233 176 -232
rect 172 -235 173 -233
rect 175 -235 176 -233
rect 178 -235 194 -232
rect 196 -234 197 -232
rect 199 -234 200 -232
rect 196 -235 200 -234
rect 222 -273 227 -272
rect 222 -275 223 -273
rect 226 -275 227 -273
rect 229 -275 231 -272
rect 234 -275 235 -272
rect 172 -279 176 -278
rect 172 -281 173 -279
rect 175 -281 176 -279
rect 178 -281 194 -278
rect 196 -280 197 -278
rect 199 -280 200 -278
rect 196 -281 200 -280
rect 222 -332 227 -331
rect 222 -334 223 -332
rect 226 -334 227 -332
rect 229 -334 231 -331
rect 234 -334 235 -331
rect 172 -338 176 -337
rect 172 -340 173 -338
rect 175 -340 176 -338
rect 178 -340 194 -337
rect 196 -339 197 -337
rect 199 -339 200 -337
rect 196 -340 200 -339
<< pdiffusion >>
rect 222 63 223 66
rect 226 63 227 66
rect 172 61 176 62
rect 172 59 173 61
rect 175 59 176 61
rect 172 57 176 59
rect 178 60 185 62
rect 178 58 179 60
rect 181 58 185 60
rect 178 57 185 58
rect 189 61 194 62
rect 189 59 190 61
rect 192 59 194 61
rect 189 57 194 59
rect 196 61 200 62
rect 196 59 197 61
rect 199 59 200 61
rect 222 60 227 63
rect 229 65 235 66
rect 229 62 231 65
rect 234 62 235 65
rect 229 60 235 62
rect 196 57 200 59
rect 222 8 223 11
rect 226 8 227 11
rect 172 6 176 7
rect 172 4 173 6
rect 175 4 176 6
rect 172 2 176 4
rect 178 5 185 7
rect 178 3 179 5
rect 181 3 185 5
rect 178 2 185 3
rect 189 6 194 7
rect 189 4 190 6
rect 192 4 194 6
rect 189 2 194 4
rect 196 6 200 7
rect 196 4 197 6
rect 199 4 200 6
rect 222 5 227 8
rect 229 10 235 11
rect 229 7 231 10
rect 234 7 235 10
rect 229 5 235 7
rect 196 2 200 4
rect 108 -22 113 -21
rect 108 -24 109 -22
rect 111 -24 113 -22
rect 108 -26 113 -24
rect 115 -26 123 -21
rect 125 -23 128 -21
rect 125 -25 126 -23
rect 125 -26 128 -25
rect 133 -22 137 -21
rect 133 -24 134 -22
rect 136 -24 137 -22
rect 133 -26 137 -24
rect 139 -23 143 -21
rect 139 -25 140 -23
rect 142 -25 143 -23
rect 139 -26 143 -25
rect 222 -38 223 -35
rect 226 -38 227 -35
rect 172 -40 176 -39
rect 172 -42 173 -40
rect 175 -42 176 -40
rect 172 -44 176 -42
rect 178 -41 185 -39
rect 178 -43 179 -41
rect 181 -43 185 -41
rect 178 -44 185 -43
rect 189 -40 194 -39
rect 189 -42 190 -40
rect 192 -42 194 -40
rect 189 -44 194 -42
rect 196 -40 200 -39
rect 196 -42 197 -40
rect 199 -42 200 -40
rect 222 -41 227 -38
rect 229 -36 235 -35
rect 229 -39 231 -36
rect 234 -39 235 -36
rect 229 -41 235 -39
rect 196 -44 200 -42
rect 222 -97 223 -94
rect 226 -97 227 -94
rect 172 -99 176 -98
rect 172 -101 173 -99
rect 175 -101 176 -99
rect 172 -103 176 -101
rect 178 -100 185 -98
rect 178 -102 179 -100
rect 181 -102 185 -100
rect 178 -103 185 -102
rect 189 -99 194 -98
rect 189 -101 190 -99
rect 192 -101 194 -99
rect 189 -103 194 -101
rect 196 -99 200 -98
rect 196 -101 197 -99
rect 199 -101 200 -99
rect 222 -100 227 -97
rect 229 -95 235 -94
rect 229 -98 231 -95
rect 234 -98 235 -95
rect 229 -100 235 -98
rect 196 -103 200 -101
rect 222 -160 223 -157
rect 226 -160 227 -157
rect 172 -162 176 -161
rect 172 -164 173 -162
rect 175 -164 176 -162
rect 172 -166 176 -164
rect 178 -163 185 -161
rect 178 -165 179 -163
rect 181 -165 185 -163
rect 178 -166 185 -165
rect 189 -162 194 -161
rect 189 -164 190 -162
rect 192 -164 194 -162
rect 189 -166 194 -164
rect 196 -162 200 -161
rect 196 -164 197 -162
rect 199 -164 200 -162
rect 222 -163 227 -160
rect 229 -158 235 -157
rect 229 -161 231 -158
rect 234 -161 235 -158
rect 229 -163 235 -161
rect 196 -166 200 -164
rect 222 -215 223 -212
rect 226 -215 227 -212
rect 172 -217 176 -216
rect 172 -219 173 -217
rect 175 -219 176 -217
rect 172 -221 176 -219
rect 178 -218 185 -216
rect 178 -220 179 -218
rect 181 -220 185 -218
rect 178 -221 185 -220
rect 189 -217 194 -216
rect 189 -219 190 -217
rect 192 -219 194 -217
rect 189 -221 194 -219
rect 196 -217 200 -216
rect 196 -219 197 -217
rect 199 -219 200 -217
rect 222 -218 227 -215
rect 229 -213 235 -212
rect 229 -216 231 -213
rect 234 -216 235 -213
rect 229 -218 235 -216
rect 196 -221 200 -219
rect 222 -261 223 -258
rect 226 -261 227 -258
rect 172 -263 176 -262
rect 172 -265 173 -263
rect 175 -265 176 -263
rect 172 -267 176 -265
rect 178 -264 185 -262
rect 178 -266 179 -264
rect 181 -266 185 -264
rect 178 -267 185 -266
rect 189 -263 194 -262
rect 189 -265 190 -263
rect 192 -265 194 -263
rect 189 -267 194 -265
rect 196 -263 200 -262
rect 196 -265 197 -263
rect 199 -265 200 -263
rect 222 -264 227 -261
rect 229 -259 235 -258
rect 229 -262 231 -259
rect 234 -262 235 -259
rect 229 -264 235 -262
rect 196 -267 200 -265
rect 222 -320 223 -317
rect 226 -320 227 -317
rect 172 -322 176 -321
rect 172 -324 173 -322
rect 175 -324 176 -322
rect 172 -326 176 -324
rect 178 -323 185 -321
rect 178 -325 179 -323
rect 181 -325 185 -323
rect 178 -326 185 -325
rect 189 -322 194 -321
rect 189 -324 190 -322
rect 192 -324 194 -322
rect 189 -326 194 -324
rect 196 -322 200 -321
rect 196 -324 197 -322
rect 199 -324 200 -322
rect 222 -323 227 -320
rect 229 -318 235 -317
rect 229 -321 231 -318
rect 234 -321 235 -318
rect 229 -323 235 -321
rect 196 -326 200 -324
<< ndcontact >>
rect 223 48 226 51
rect 231 49 234 52
rect 173 43 175 45
rect 197 44 199 46
rect 223 -7 226 -4
rect 231 -6 234 -3
rect 173 -12 175 -10
rect 197 -11 199 -9
rect 110 -38 112 -36
rect 116 -38 118 -36
rect 120 -38 122 -36
rect 126 -38 128 -36
rect 134 -38 136 -36
rect 140 -38 142 -36
rect 223 -53 226 -50
rect 231 -52 234 -49
rect 173 -58 175 -56
rect 197 -57 199 -55
rect 223 -112 226 -109
rect 231 -111 234 -108
rect 173 -117 175 -115
rect 197 -116 199 -114
rect 223 -175 226 -172
rect 231 -174 234 -171
rect 173 -180 175 -178
rect 197 -179 199 -177
rect 223 -230 226 -227
rect 231 -229 234 -226
rect 173 -235 175 -233
rect 197 -234 199 -232
rect 223 -276 226 -273
rect 231 -275 234 -272
rect 173 -281 175 -279
rect 197 -280 199 -278
rect 223 -335 226 -332
rect 231 -334 234 -331
rect 173 -340 175 -338
rect 197 -339 199 -337
<< pdcontact >>
rect 223 63 226 66
rect 173 59 175 61
rect 179 58 181 60
rect 190 59 192 61
rect 197 59 199 61
rect 231 62 234 65
rect 223 8 226 11
rect 173 4 175 6
rect 179 3 181 5
rect 190 4 192 6
rect 197 4 199 6
rect 231 7 234 10
rect 109 -24 111 -22
rect 126 -25 128 -23
rect 134 -24 136 -22
rect 140 -25 142 -23
rect 223 -38 226 -35
rect 173 -42 175 -40
rect 179 -43 181 -41
rect 190 -42 192 -40
rect 197 -42 199 -40
rect 231 -39 234 -36
rect 223 -97 226 -94
rect 173 -101 175 -99
rect 179 -102 181 -100
rect 190 -101 192 -99
rect 197 -101 199 -99
rect 231 -98 234 -95
rect 223 -160 226 -157
rect 173 -164 175 -162
rect 179 -165 181 -163
rect 190 -164 192 -162
rect 197 -164 199 -162
rect 231 -161 234 -158
rect 223 -215 226 -212
rect 173 -219 175 -217
rect 179 -220 181 -218
rect 190 -219 192 -217
rect 197 -219 199 -217
rect 231 -216 234 -213
rect 223 -261 226 -258
rect 173 -265 175 -263
rect 179 -266 181 -264
rect 190 -265 192 -263
rect 197 -265 199 -263
rect 231 -262 234 -259
rect 223 -320 226 -317
rect 173 -324 175 -322
rect 179 -325 181 -323
rect 190 -324 192 -322
rect 197 -324 199 -322
rect 231 -321 234 -318
<< polysilicon >>
rect 227 66 229 79
rect 176 62 178 65
rect 194 62 196 65
rect 176 50 178 57
rect 157 48 178 50
rect 157 -5 159 48
rect 176 46 178 48
rect 194 46 196 57
rect 227 56 229 60
rect 228 53 229 56
rect 227 52 229 53
rect 227 47 229 49
rect 176 42 178 43
rect 194 42 196 43
rect 227 11 229 24
rect 176 7 178 10
rect 194 7 196 10
rect 176 -5 178 2
rect 157 -7 178 -5
rect 113 -21 115 -19
rect 123 -21 125 -19
rect 137 -21 139 -19
rect 113 -36 115 -26
rect 123 -36 125 -26
rect 137 -31 139 -26
rect 157 -31 159 -7
rect 176 -9 178 -7
rect 194 -9 196 2
rect 227 1 229 5
rect 228 -2 229 1
rect 227 -3 229 -2
rect 227 -8 229 -6
rect 176 -13 178 -12
rect 194 -13 196 -12
rect 138 -33 139 -31
rect 147 -33 159 -31
rect 137 -36 139 -33
rect 113 -40 115 -39
rect 123 -40 125 -39
rect 137 -40 139 -39
rect 157 -52 159 -33
rect 227 -35 229 -22
rect 176 -39 178 -36
rect 194 -39 196 -36
rect 176 -52 178 -44
rect 157 -54 178 -52
rect 157 -110 159 -54
rect 176 -55 178 -54
rect 194 -55 196 -44
rect 227 -45 229 -41
rect 228 -48 229 -45
rect 227 -49 229 -48
rect 227 -54 229 -52
rect 176 -59 178 -58
rect 194 -59 196 -58
rect 227 -94 229 -81
rect 176 -98 178 -95
rect 194 -98 196 -95
rect 176 -110 178 -103
rect 157 -112 178 -110
rect 157 -173 159 -112
rect 176 -114 178 -112
rect 194 -114 196 -103
rect 227 -104 229 -100
rect 228 -107 229 -104
rect 227 -108 229 -107
rect 227 -113 229 -111
rect 176 -118 178 -117
rect 194 -118 196 -117
rect 227 -157 229 -144
rect 176 -161 178 -158
rect 194 -161 196 -158
rect 176 -173 178 -166
rect 157 -175 178 -173
rect 157 -228 159 -175
rect 176 -177 178 -175
rect 194 -177 196 -166
rect 227 -167 229 -163
rect 228 -170 229 -167
rect 227 -171 229 -170
rect 227 -176 229 -174
rect 176 -181 178 -180
rect 194 -181 196 -180
rect 227 -212 229 -199
rect 176 -216 178 -213
rect 194 -216 196 -213
rect 176 -228 178 -221
rect 157 -230 178 -228
rect 157 -254 159 -230
rect 176 -232 178 -230
rect 194 -232 196 -221
rect 227 -222 229 -218
rect 228 -225 229 -222
rect 227 -226 229 -225
rect 227 -231 229 -229
rect 176 -236 178 -235
rect 194 -236 196 -235
rect 156 -256 159 -254
rect 157 -275 159 -256
rect 227 -258 229 -245
rect 176 -262 178 -259
rect 194 -262 196 -259
rect 176 -275 178 -267
rect 157 -277 178 -275
rect 157 -333 159 -277
rect 176 -278 178 -277
rect 194 -278 196 -267
rect 227 -268 229 -264
rect 228 -271 229 -268
rect 227 -272 229 -271
rect 227 -277 229 -275
rect 176 -282 178 -281
rect 194 -282 196 -281
rect 227 -317 229 -304
rect 176 -321 178 -318
rect 194 -321 196 -318
rect 176 -333 178 -326
rect 157 -335 178 -333
rect 176 -337 178 -335
rect 194 -337 196 -326
rect 227 -327 229 -323
rect 228 -330 229 -327
rect 227 -331 229 -330
rect 227 -336 229 -334
rect 176 -341 178 -340
rect 194 -341 196 -340
<< polycontact >>
rect 225 53 228 56
rect 225 -2 228 1
rect 137 -33 138 -31
rect 142 -33 147 -31
rect 225 -48 228 -45
rect 225 -107 228 -104
rect 225 -170 228 -167
rect 225 -225 228 -222
rect 225 -271 228 -268
rect 225 -330 228 -327
<< metal1 >>
rect 223 72 249 74
rect 223 69 226 72
rect 134 67 226 69
rect 134 -16 136 67
rect 173 61 175 67
rect 190 61 192 67
rect 223 66 226 67
rect 179 52 181 58
rect 197 52 199 59
rect 231 57 234 62
rect 215 53 225 56
rect 231 54 237 57
rect 215 52 217 53
rect 179 50 217 52
rect 231 52 234 54
rect 197 46 199 50
rect 223 45 226 48
rect 173 41 175 43
rect 223 43 234 45
rect 223 41 227 43
rect 161 39 227 41
rect 161 -14 163 39
rect 247 19 249 72
rect 223 17 249 19
rect 223 14 226 17
rect 173 12 226 14
rect 173 6 175 12
rect 190 6 192 12
rect 223 11 226 12
rect 179 -3 181 3
rect 197 -3 199 4
rect 231 2 234 7
rect 215 -2 225 1
rect 231 -1 237 2
rect 215 -3 217 -2
rect 179 -5 217 -3
rect 231 -3 234 -1
rect 197 -9 199 -5
rect 223 -10 226 -7
rect 173 -14 175 -12
rect 223 -12 234 -10
rect 223 -14 227 -12
rect 161 -16 227 -14
rect 109 -18 139 -16
rect 109 -22 111 -18
rect 134 -22 136 -18
rect 126 -31 128 -25
rect 116 -33 137 -31
rect 116 -36 118 -33
rect 126 -36 128 -33
rect 140 -36 142 -25
rect 110 -41 112 -38
rect 120 -41 122 -38
rect 134 -41 136 -38
rect 161 -41 163 -16
rect 247 -27 249 17
rect 223 -29 249 -27
rect 223 -32 226 -29
rect 108 -43 163 -41
rect 173 -34 226 -32
rect 173 -40 175 -34
rect 190 -40 192 -34
rect 223 -35 226 -34
rect 161 -60 163 -43
rect 179 -49 181 -43
rect 197 -49 199 -42
rect 231 -44 234 -39
rect 215 -48 225 -45
rect 231 -47 237 -44
rect 215 -49 217 -48
rect 179 -51 217 -49
rect 231 -49 234 -47
rect 197 -55 199 -51
rect 223 -56 226 -53
rect 173 -60 175 -58
rect 223 -58 234 -56
rect 223 -60 227 -58
rect 161 -62 227 -60
rect 161 -119 163 -62
rect 247 -86 249 -29
rect 223 -88 249 -86
rect 223 -91 226 -88
rect 173 -93 226 -91
rect 173 -99 175 -93
rect 190 -99 192 -93
rect 223 -94 226 -93
rect 179 -108 181 -102
rect 197 -108 199 -101
rect 231 -103 234 -98
rect 215 -107 225 -104
rect 231 -106 237 -103
rect 215 -108 217 -107
rect 179 -110 217 -108
rect 231 -108 234 -106
rect 197 -114 199 -110
rect 223 -115 226 -112
rect 173 -119 175 -117
rect 223 -117 234 -115
rect 223 -119 227 -117
rect 161 -121 227 -119
rect 161 -182 163 -121
rect 247 -149 249 -88
rect 223 -151 249 -149
rect 223 -154 226 -151
rect 168 -156 226 -154
rect 173 -162 175 -156
rect 190 -162 192 -156
rect 223 -157 226 -156
rect 179 -171 181 -165
rect 197 -171 199 -164
rect 231 -166 234 -161
rect 215 -170 225 -167
rect 231 -169 237 -166
rect 215 -171 217 -170
rect 179 -173 217 -171
rect 231 -171 234 -169
rect 197 -177 199 -173
rect 223 -178 226 -175
rect 173 -182 175 -180
rect 223 -180 234 -178
rect 223 -182 227 -180
rect 161 -184 227 -182
rect 161 -237 163 -184
rect 247 -204 249 -151
rect 223 -206 249 -204
rect 223 -209 226 -206
rect 173 -211 226 -209
rect 173 -217 175 -211
rect 190 -217 192 -211
rect 223 -212 226 -211
rect 179 -226 181 -220
rect 197 -226 199 -219
rect 231 -221 234 -216
rect 215 -225 225 -222
rect 231 -224 237 -221
rect 215 -226 217 -225
rect 179 -228 217 -226
rect 231 -226 234 -224
rect 197 -232 199 -228
rect 223 -233 226 -230
rect 173 -237 175 -235
rect 223 -235 234 -233
rect 223 -237 227 -235
rect 161 -239 227 -237
rect 161 -264 163 -239
rect 247 -250 249 -206
rect 223 -252 249 -250
rect 223 -255 226 -252
rect 156 -266 163 -264
rect 173 -257 226 -255
rect 173 -263 175 -257
rect 190 -263 192 -257
rect 223 -258 226 -257
rect 161 -283 163 -266
rect 179 -272 181 -266
rect 197 -272 199 -265
rect 231 -267 234 -262
rect 215 -271 225 -268
rect 231 -270 237 -267
rect 215 -272 217 -271
rect 179 -274 217 -272
rect 231 -272 234 -270
rect 197 -278 199 -274
rect 223 -279 226 -276
rect 173 -283 175 -281
rect 223 -281 234 -279
rect 223 -283 227 -281
rect 161 -285 227 -283
rect 161 -342 163 -285
rect 247 -309 249 -252
rect 223 -311 249 -309
rect 223 -314 226 -311
rect 173 -316 226 -314
rect 173 -322 175 -316
rect 190 -322 192 -316
rect 223 -317 226 -316
rect 179 -331 181 -325
rect 197 -331 199 -324
rect 231 -326 234 -321
rect 215 -330 225 -327
rect 231 -329 237 -326
rect 215 -331 217 -330
rect 179 -333 217 -331
rect 231 -331 234 -329
rect 197 -337 199 -333
rect 223 -338 226 -335
rect 173 -342 175 -340
rect 223 -340 234 -338
rect 223 -342 227 -340
rect 161 -344 227 -342
<< labels >>
rlabel polysilicon 114 -32 114 -32 1 D0
rlabel polysilicon 124 -35 124 -35 1 D1
rlabel polysilicon 152 -32 152 -32 1 D
rlabel metal1 131 -42 131 -42 1 gnd
rlabel metal1 124 -17 124 -17 1 vdd
rlabel polysilicon 195 -53 195 -53 1 a1
rlabel polysilicon 195 -7 195 -7 1 a2
rlabel polysilicon 195 49 195 49 1 a3
rlabel metal1 234 56 234 56 1 adsub_a3
rlabel metal1 235 0 235 0 1 adsub_a2
rlabel metal1 235 -46 235 -46 1 adsub_a1
rlabel metal1 235 -105 235 -105 1 adsub_a0
rlabel polysilicon 195 -112 195 -112 1 a0
rlabel polysilicon 195 -174 195 -174 1 b3
rlabel metal1 235 -168 235 -168 1 adsub_b3
rlabel polysilicon 195 -230 195 -230 1 b2
rlabel metal1 235 -222 235 -222 1 adsub_b2
rlabel polysilicon 195 -276 195 -276 1 b1
rlabel metal1 234 -268 234 -268 1 adsub_b1
rlabel polysilicon 195 -335 195 -335 1 b0
rlabel metal1 235 -327 235 -327 1 adsub_b0
<< end >>
