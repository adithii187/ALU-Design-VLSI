magic
tech scmos
timestamp 1700473287
<< error_p >>
rect -167 334 -166 335
rect -166 333 -165 334
<< nwell >>
rect -756 108 -648 783
rect 54 108 162 783
rect 936 108 1044 783
rect 594 -81 783 -27
rect -432 -144 -243 -90
rect -900 -297 -576 -207
rect -432 -252 -279 -144
rect 126 -234 450 -144
rect 594 -189 747 -81
rect 594 -198 657 -189
rect 675 -198 747 -189
rect -432 -261 -369 -252
rect -351 -261 -279 -252
rect -216 -648 135 -531
<< ntransistor >>
rect -981 702 -927 720
rect -171 702 -117 720
rect -981 531 -927 549
rect -981 333 -927 351
rect -981 171 -927 189
rect 711 702 765 720
rect -171 531 -117 549
rect -171 334 -117 351
rect -166 333 -117 334
rect -171 171 -117 189
rect 711 531 765 549
rect 711 333 765 351
rect 711 171 765 189
rect -369 -342 -351 -315
rect -828 -396 -810 -369
rect -666 -396 -648 -369
rect 198 -333 216 -306
rect 360 -333 378 -306
rect 657 -279 675 -252
rect -153 -747 -135 -720
rect -63 -747 -45 -720
rect 63 -747 81 -720
<< ptransistor >>
rect -729 702 -666 720
rect 81 702 144 720
rect -729 531 -666 549
rect -729 333 -666 351
rect -729 171 -666 189
rect 963 702 1026 720
rect 81 531 144 549
rect 81 333 144 351
rect 81 171 144 189
rect 963 531 1026 549
rect 963 333 1026 351
rect 963 171 1026 189
rect -828 -270 -810 -225
rect -666 -270 -648 -225
rect -369 -243 -351 -189
rect 198 -207 216 -162
rect 360 -207 378 -162
rect 657 -180 675 -126
rect -153 -630 -135 -585
rect -63 -630 -45 -585
rect 63 -630 81 -585
<< ndiffusion >>
rect -981 765 -927 774
rect -981 729 -972 765
rect -936 729 -927 765
rect -981 720 -927 729
rect -981 693 -927 702
rect -981 657 -972 693
rect -936 657 -927 693
rect -981 648 -927 657
rect -981 594 -927 603
rect -981 558 -972 594
rect -936 558 -927 594
rect -981 549 -927 558
rect -171 765 -117 774
rect -171 729 -162 765
rect -126 729 -117 765
rect -171 720 -117 729
rect -981 522 -927 531
rect -981 486 -972 522
rect -936 486 -927 522
rect -981 477 -927 486
rect -981 405 -927 414
rect -981 369 -972 405
rect -936 369 -927 405
rect -981 351 -927 369
rect -981 324 -927 333
rect -981 288 -972 324
rect -936 288 -927 324
rect -981 279 -927 288
rect -981 243 -927 252
rect -981 207 -972 243
rect -936 207 -927 243
rect -981 189 -927 207
rect -981 162 -927 171
rect -981 126 -972 162
rect -936 126 -927 162
rect -981 117 -927 126
rect -171 693 -117 702
rect -171 657 -162 693
rect -126 657 -117 693
rect -171 648 -117 657
rect -171 594 -117 603
rect -171 558 -162 594
rect -126 558 -117 594
rect -171 549 -117 558
rect 711 765 765 774
rect 711 729 720 765
rect 756 729 765 765
rect 711 720 765 729
rect -171 522 -117 531
rect -171 486 -162 522
rect -126 486 -117 522
rect -171 477 -117 486
rect -171 405 -117 414
rect -171 369 -162 405
rect -126 369 -117 405
rect -171 351 -117 369
rect -171 333 -166 334
rect -171 324 -117 333
rect -171 288 -162 324
rect -126 288 -117 324
rect -171 279 -117 288
rect -171 243 -117 252
rect -171 207 -162 243
rect -126 207 -117 243
rect -171 189 -117 207
rect -171 162 -117 171
rect -171 126 -162 162
rect -126 126 -117 162
rect -171 117 -117 126
rect 711 693 765 702
rect 711 657 720 693
rect 756 657 765 693
rect 711 648 765 657
rect 711 594 765 603
rect 711 558 720 594
rect 756 558 765 594
rect 711 549 765 558
rect 711 522 765 531
rect 711 486 720 522
rect 756 486 765 522
rect 711 477 765 486
rect 711 405 765 414
rect 711 369 720 405
rect 756 369 765 405
rect 711 351 765 369
rect 711 324 765 333
rect 711 288 720 324
rect 756 288 765 324
rect 711 279 765 288
rect 711 243 765 252
rect 711 207 720 243
rect 756 207 765 243
rect 711 189 765 207
rect 711 162 765 171
rect 711 126 720 162
rect 756 126 765 162
rect 711 117 765 126
rect -414 -324 -369 -315
rect -414 -342 -405 -324
rect -378 -342 -369 -324
rect -351 -342 -333 -315
rect -306 -342 -297 -315
rect -864 -378 -828 -369
rect -864 -396 -855 -378
rect -837 -396 -828 -378
rect -810 -396 -666 -369
rect -648 -387 -639 -369
rect -621 -387 -612 -369
rect -648 -396 -612 -387
rect 162 -315 198 -306
rect 162 -333 171 -315
rect 189 -333 198 -315
rect 216 -333 360 -306
rect 378 -324 387 -306
rect 405 -324 414 -306
rect 378 -333 414 -324
rect 612 -261 657 -252
rect 612 -279 621 -261
rect 648 -279 657 -261
rect 675 -279 693 -252
rect 720 -279 729 -252
rect -189 -738 -180 -720
rect -162 -738 -153 -720
rect -189 -747 -153 -738
rect -135 -738 -126 -720
rect -135 -747 -108 -738
rect -99 -738 -90 -720
rect -72 -738 -63 -720
rect -99 -747 -63 -738
rect -45 -738 -36 -720
rect -45 -747 -18 -738
rect 27 -738 36 -720
rect 54 -738 63 -720
rect 27 -747 63 -738
rect 81 -738 90 -720
rect 108 -738 117 -720
rect 81 -747 117 -738
<< pdiffusion >>
rect -729 765 -666 774
rect -729 729 -720 765
rect -684 729 -666 765
rect -729 720 -666 729
rect -729 693 -666 702
rect -729 657 -720 693
rect -684 657 -666 693
rect -729 648 -666 657
rect -729 594 -666 603
rect -729 558 -720 594
rect -684 558 -666 594
rect -729 549 -666 558
rect 81 765 144 774
rect 81 729 90 765
rect 126 729 144 765
rect 81 720 144 729
rect -729 522 -666 531
rect -729 486 -720 522
rect -684 486 -666 522
rect -729 477 -666 486
rect -729 405 -666 414
rect -729 369 -720 405
rect -684 369 -666 405
rect -729 351 -666 369
rect -729 324 -666 333
rect -729 288 -720 324
rect -684 288 -666 324
rect -729 279 -666 288
rect -729 243 -666 252
rect -729 207 -720 243
rect -684 207 -666 243
rect -729 189 -666 207
rect -729 162 -666 171
rect -729 126 -720 162
rect -684 126 -666 162
rect -729 117 -666 126
rect 81 693 144 702
rect 81 657 90 693
rect 126 657 144 693
rect 81 648 144 657
rect 81 594 144 603
rect 81 558 90 594
rect 126 558 144 594
rect 81 549 144 558
rect 963 765 1026 774
rect 963 729 972 765
rect 1008 729 1026 765
rect 963 720 1026 729
rect 81 522 144 531
rect 81 486 90 522
rect 126 486 144 522
rect 81 477 144 486
rect 81 405 144 414
rect 81 369 90 405
rect 126 369 144 405
rect 81 351 144 369
rect 81 324 144 333
rect 81 288 90 324
rect 126 288 144 324
rect 81 279 144 288
rect 81 243 144 252
rect 81 207 90 243
rect 126 207 144 243
rect 81 189 144 207
rect 81 162 144 171
rect 81 126 90 162
rect 126 126 144 162
rect 81 117 144 126
rect 963 693 1026 702
rect 963 657 972 693
rect 1008 657 1026 693
rect 963 648 1026 657
rect 963 594 1026 603
rect 963 558 972 594
rect 1008 558 1026 594
rect 963 549 1026 558
rect 963 522 1026 531
rect 963 486 972 522
rect 1008 486 1026 522
rect 963 477 1026 486
rect 963 405 1026 414
rect 963 369 972 405
rect 1008 369 1026 405
rect 963 351 1026 369
rect 963 324 1026 333
rect 963 288 972 324
rect 1008 288 1026 324
rect 963 279 1026 288
rect 963 243 1026 252
rect 963 207 972 243
rect 1008 207 1026 243
rect 963 189 1026 207
rect 963 162 1026 171
rect 963 126 972 162
rect 1008 126 1026 162
rect 963 117 1026 126
rect -864 -234 -828 -225
rect -864 -252 -855 -234
rect -837 -252 -828 -234
rect -864 -270 -828 -252
rect -810 -243 -747 -225
rect -810 -261 -801 -243
rect -783 -261 -747 -243
rect -810 -270 -747 -261
rect -711 -234 -666 -225
rect -711 -252 -702 -234
rect -684 -252 -666 -234
rect -711 -270 -666 -252
rect -648 -234 -612 -225
rect -648 -252 -639 -234
rect -621 -252 -612 -234
rect -648 -270 -612 -252
rect -414 -216 -405 -189
rect -378 -216 -369 -189
rect -414 -243 -369 -216
rect -351 -198 -297 -189
rect -351 -225 -333 -198
rect -306 -225 -297 -198
rect -351 -243 -297 -225
rect 162 -171 198 -162
rect 162 -189 171 -171
rect 189 -189 198 -171
rect 162 -207 198 -189
rect 216 -180 279 -162
rect 216 -198 225 -180
rect 243 -198 279 -180
rect 216 -207 279 -198
rect 315 -171 360 -162
rect 315 -189 324 -171
rect 342 -189 360 -171
rect 315 -207 360 -189
rect 378 -171 414 -162
rect 378 -189 387 -171
rect 405 -189 414 -171
rect 378 -207 414 -189
rect 612 -153 621 -126
rect 648 -153 657 -126
rect 612 -180 657 -153
rect 675 -135 729 -126
rect 675 -162 693 -135
rect 720 -162 729 -135
rect 675 -180 729 -162
rect -198 -594 -153 -585
rect -198 -612 -189 -594
rect -171 -612 -153 -594
rect -198 -630 -153 -612
rect -135 -630 -63 -585
rect -45 -603 -18 -585
rect -45 -621 -36 -603
rect -45 -630 -18 -621
rect 27 -594 63 -585
rect 27 -612 36 -594
rect 54 -612 63 -594
rect 27 -630 63 -612
rect 81 -603 117 -585
rect 81 -621 90 -603
rect 108 -621 117 -603
rect 81 -630 117 -621
<< ndcontact >>
rect -972 729 -936 765
rect -972 657 -936 693
rect -972 558 -936 594
rect -162 729 -126 765
rect -972 486 -936 522
rect -972 369 -936 405
rect -972 288 -936 324
rect -972 207 -936 243
rect -972 126 -936 162
rect -162 657 -126 693
rect -162 558 -126 594
rect 720 729 756 765
rect -162 486 -126 522
rect -162 369 -126 405
rect -162 288 -126 324
rect -162 207 -126 243
rect -162 126 -126 162
rect 720 657 756 693
rect 720 558 756 594
rect 720 486 756 522
rect 720 369 756 405
rect 720 288 756 324
rect 720 207 756 243
rect 720 126 756 162
rect -405 -351 -378 -324
rect -333 -342 -306 -315
rect -855 -396 -837 -378
rect -639 -387 -621 -369
rect 171 -333 189 -315
rect 387 -324 405 -306
rect 621 -288 648 -261
rect 693 -279 720 -252
rect -180 -738 -162 -720
rect -126 -738 -108 -720
rect -90 -738 -72 -720
rect -36 -738 -18 -720
rect 36 -738 54 -720
rect 90 -738 108 -720
<< pdcontact >>
rect -720 729 -684 765
rect -720 657 -684 693
rect -720 558 -684 594
rect 90 729 126 765
rect -720 486 -684 522
rect -720 369 -684 405
rect -720 288 -684 324
rect -720 207 -684 243
rect -720 126 -684 162
rect 90 657 126 693
rect 90 558 126 594
rect 972 729 1008 765
rect 90 486 126 522
rect 90 369 126 405
rect 90 288 126 324
rect 90 207 126 243
rect 90 126 126 162
rect 972 657 1008 693
rect 972 558 1008 594
rect 972 486 1008 522
rect 972 369 1008 405
rect 972 288 1008 324
rect 972 207 1008 243
rect 972 126 1008 162
rect -855 -252 -837 -234
rect -801 -261 -783 -243
rect -702 -252 -684 -234
rect -639 -252 -621 -234
rect -405 -216 -378 -189
rect -333 -225 -306 -198
rect 171 -189 189 -171
rect 225 -198 243 -180
rect 324 -189 342 -171
rect 387 -189 405 -171
rect 621 -153 648 -126
rect 693 -162 720 -135
rect -189 -612 -171 -594
rect -36 -621 -18 -603
rect 36 -612 54 -594
rect 90 -621 108 -603
<< psubstratepcontact >>
rect -1098 333 -1062 369
rect -1098 243 -1062 279
rect -288 333 -252 369
rect -288 243 -252 279
rect 594 333 630 369
rect 594 243 630 279
<< nsubstratencontact >>
rect -603 333 -567 369
rect -603 243 -567 279
rect 207 333 243 369
rect 207 243 243 279
rect 1089 333 1125 369
rect 1089 243 1125 279
<< polysilicon >>
rect -1035 810 -594 828
rect -1035 720 -1017 810
rect -1188 702 -981 720
rect -927 702 -918 720
rect -900 702 -729 720
rect -666 702 -639 720
rect -1188 63 -1170 702
rect -900 549 -882 702
rect -612 549 -594 810
rect -225 810 216 828
rect -225 720 -207 810
rect -378 702 -171 720
rect -117 702 -108 720
rect -90 702 81 720
rect 144 702 171 720
rect -549 603 -450 621
rect -1143 531 -981 549
rect -927 531 -882 549
rect -765 531 -729 549
rect -666 531 -594 549
rect -1143 189 -1125 531
rect -855 351 -819 378
rect -1044 333 -981 351
rect -927 333 -729 351
rect -666 333 -621 351
rect -468 342 -450 603
rect -522 324 -450 342
rect -855 189 -819 234
rect -1143 171 -981 189
rect -927 171 -729 189
rect -666 171 -621 189
rect -1188 45 -819 63
rect -522 45 -504 324
rect -468 315 -450 324
rect -443 297 -441 315
rect -378 63 -360 702
rect -90 549 -72 702
rect 198 549 216 810
rect 657 810 1098 828
rect 657 720 675 810
rect 504 702 711 720
rect 765 702 774 720
rect 792 702 963 720
rect 1026 702 1053 720
rect 261 603 387 621
rect -333 531 -171 549
rect -117 531 -72 549
rect 45 531 81 549
rect 144 531 216 549
rect -333 315 -315 531
rect -45 351 -9 378
rect -234 334 -171 351
rect -117 333 81 351
rect 144 333 189 351
rect -333 297 -312 315
rect -333 189 -315 297
rect -36 270 -18 333
rect 369 315 387 603
rect 369 297 414 315
rect -185 261 -18 270
rect -45 189 -9 234
rect -333 171 -171 189
rect -117 171 81 189
rect 144 171 189 189
rect -378 45 -9 63
rect -657 27 -504 45
rect -657 -81 -639 27
rect 18 -36 36 171
rect 369 -18 387 297
rect 438 297 450 315
rect 504 63 522 702
rect 792 549 810 702
rect 1080 549 1098 810
rect 1143 594 1224 630
rect 549 531 711 549
rect 765 531 810 549
rect 927 531 963 549
rect 1026 531 1098 549
rect 549 337 567 531
rect 549 285 568 337
rect 837 351 873 378
rect 648 333 711 351
rect 765 333 963 351
rect 1026 333 1071 351
rect 549 189 567 285
rect 846 270 864 333
rect 700 261 864 270
rect 837 189 873 234
rect 549 171 711 189
rect 765 171 963 189
rect 1026 171 1071 189
rect 504 45 873 63
rect 900 27 918 171
rect -927 -99 -639 -81
rect -549 -54 36 -36
rect 99 -36 387 -18
rect 477 9 918 27
rect -927 -333 -909 -99
rect -828 -225 -810 -198
rect -666 -225 -648 -198
rect -828 -333 -810 -270
rect -927 -351 -810 -333
rect -828 -369 -810 -351
rect -666 -342 -648 -270
rect -549 -342 -531 -54
rect -369 -189 -351 -72
rect -369 -279 -351 -243
rect -360 -306 -351 -279
rect -369 -315 -351 -306
rect -666 -360 -531 -342
rect -369 -360 -351 -342
rect -666 -369 -648 -360
rect -828 -405 -810 -396
rect -666 -405 -648 -396
rect -270 -675 -252 -270
rect -108 -540 -90 -135
rect -27 -378 -9 -90
rect 99 -270 117 -36
rect 198 -162 216 -135
rect 360 -162 378 -135
rect 198 -270 216 -207
rect 99 -288 216 -270
rect 198 -306 216 -288
rect 360 -279 378 -207
rect 477 -279 495 9
rect 360 -297 495 -279
rect 360 -306 378 -297
rect 198 -342 216 -333
rect 360 -342 378 -333
rect 513 -351 531 -18
rect 657 -126 675 -9
rect 657 -216 675 -180
rect 666 -243 675 -216
rect 756 -234 792 -207
rect 657 -252 675 -243
rect 657 -297 675 -279
rect 774 -423 792 -234
rect 0 -441 792 -423
rect -153 -585 -135 -567
rect -63 -585 -45 -567
rect -153 -675 -135 -630
rect -270 -693 -135 -675
rect -153 -720 -135 -693
rect -63 -702 -45 -630
rect 0 -702 18 -441
rect 63 -585 81 -567
rect -63 -711 18 -702
rect 63 -675 81 -630
rect 72 -693 81 -675
rect -63 -720 -45 -711
rect 63 -720 81 -693
rect -153 -756 -135 -747
rect -63 -756 -45 -747
rect 63 -756 81 -747
<< polycontact >>
rect -585 603 -549 621
rect -855 378 -819 414
rect -855 63 -819 99
rect -468 297 -443 315
rect 225 603 261 621
rect -45 378 -9 414
rect -214 254 -185 286
rect -45 63 -9 99
rect 414 293 438 322
rect 1107 585 1143 630
rect 837 378 873 414
rect 674 253 700 279
rect 837 63 873 99
rect -36 -90 -9 -72
rect -108 -135 -90 -117
rect -387 -306 -360 -279
rect -306 -297 -270 -270
rect 513 -18 531 0
rect 639 -243 666 -216
rect 720 -234 756 -207
rect 513 -369 531 -351
rect -27 -396 -9 -378
rect -108 -558 -90 -540
rect 63 -693 72 -675
<< metal1 >>
rect -936 729 -720 765
rect -684 729 -504 765
rect -126 729 90 765
rect 126 729 306 765
rect 756 729 972 765
rect 1008 729 1188 765
rect -936 657 -720 693
rect -684 657 -549 693
rect -585 621 -549 657
rect -1098 558 -972 594
rect -936 558 -720 594
rect -1098 459 -1062 558
rect -585 522 -549 603
rect -936 486 -720 522
rect -684 486 -549 522
rect -540 459 -504 729
rect -126 657 90 693
rect 126 657 261 693
rect 225 621 261 657
rect -1098 423 -873 459
rect -1098 369 -972 405
rect -1098 306 -1062 333
rect -909 324 -873 423
rect -855 423 -504 459
rect -288 558 -162 594
rect -126 558 90 594
rect -288 459 -252 558
rect 225 522 261 603
rect -126 486 90 522
rect 126 486 261 522
rect 270 459 306 729
rect 756 657 972 693
rect 1008 657 1143 693
rect 1107 630 1143 657
rect -288 423 -63 459
rect -855 414 -819 423
rect -684 369 -567 405
rect -1251 288 -1062 306
rect -936 288 -720 324
rect -603 306 -567 333
rect -288 369 -162 405
rect -447 315 -391 321
rect -603 288 -477 306
rect -443 298 -391 315
rect -1251 -414 -1233 288
rect -1098 279 -1062 288
rect -603 279 -567 288
rect -1098 207 -972 243
rect -684 207 -567 243
rect -936 126 -720 162
rect -855 99 -819 126
rect -495 -162 -477 288
rect -288 279 -252 333
rect -99 324 -63 423
rect -45 423 306 459
rect 594 558 720 594
rect 756 558 972 594
rect 594 459 630 558
rect 1107 522 1143 585
rect 756 486 972 522
rect 1008 486 1143 522
rect 1152 459 1188 729
rect 594 423 819 459
rect -45 414 -9 423
rect 126 369 243 405
rect -214 286 -195 294
rect -126 288 90 324
rect 207 315 243 333
rect 594 369 720 405
rect 207 297 324 315
rect 207 279 243 297
rect -288 207 -162 243
rect 126 207 243 243
rect -216 -72 -198 207
rect -126 126 90 162
rect -45 99 -9 126
rect -216 -90 -36 -72
rect 306 -99 324 297
rect 438 296 467 316
rect 594 315 630 333
rect 783 324 819 423
rect 837 423 1188 459
rect 837 414 873 423
rect 1008 369 1125 405
rect 593 297 630 315
rect 594 279 630 297
rect 673 279 693 292
rect 756 288 972 324
rect 1089 315 1125 333
rect 1089 297 1170 315
rect 1089 279 1125 297
rect 673 263 674 279
rect 594 207 720 243
rect 1008 207 1125 243
rect 621 0 639 207
rect 756 126 972 162
rect 837 99 873 126
rect 531 -18 639 0
rect 1152 -54 1170 297
rect 621 -72 1170 -54
rect 621 -99 648 -72
rect 171 -117 648 -99
rect -405 -135 -108 -117
rect -90 -135 189 -117
rect -405 -162 -378 -135
rect -855 -180 -378 -162
rect -855 -234 -837 -180
rect -702 -234 -684 -180
rect -405 -189 -378 -180
rect 171 -171 189 -135
rect 324 -171 342 -117
rect 621 -126 648 -117
rect -801 -315 -783 -261
rect -639 -315 -621 -252
rect -477 -306 -387 -279
rect -477 -315 -459 -306
rect -801 -333 -459 -315
rect -333 -315 -306 -225
rect 225 -252 243 -198
rect 387 -252 405 -189
rect 549 -243 639 -216
rect 549 -252 567 -243
rect 225 -270 567 -252
rect 693 -252 720 -162
rect 387 -306 405 -270
rect -639 -369 -621 -333
rect 621 -315 648 -288
rect -405 -378 -378 -351
rect 171 -351 189 -333
rect 621 -333 720 -315
rect 621 -351 657 -333
rect 171 -369 513 -351
rect 531 -369 657 -351
rect 171 -378 189 -369
rect -855 -414 -837 -396
rect -405 -396 -27 -378
rect -9 -396 189 -378
rect -405 -414 -369 -396
rect -1251 -432 -369 -414
rect -387 -765 -369 -432
rect -189 -558 -108 -540
rect -90 -558 81 -540
rect -189 -594 -171 -558
rect 36 -594 54 -558
rect -36 -675 -18 -621
rect 90 -675 108 -621
rect -126 -693 63 -675
rect 90 -693 135 -675
rect -126 -720 -108 -693
rect -36 -720 -18 -693
rect 90 -720 108 -693
rect -180 -765 -162 -738
rect -90 -765 -72 -738
rect 36 -765 54 -738
rect -387 -783 54 -765
<< m2contact >>
rect -391 298 -362 330
rect -214 294 -185 326
rect 467 285 497 316
rect 672 292 702 323
<< metal2 >>
rect -392 298 -391 320
rect -362 298 -214 320
rect 484 316 672 317
rect 497 292 672 316
<< labels >>
rlabel polysilicon -837 207 -837 207 1 b
rlabel polysilicon -837 360 -837 360 1 m
rlabel polysilicon -27 189 -27 189 1 a
rlabel metal1 243 567 243 567 1 xor1
rlabel polysilicon 855 189 855 189 1 carry
rlabel polysilicon 1206 612 1206 612 7 sum
rlabel metal1 117 -684 117 -684 1 carry_out
rlabel metal1 -162 -774 -162 -774 1 gnd
rlabel metal1 -144 -549 -144 -549 1 vdd
rlabel polysilicon -459 603 -459 603 1 inp
rlabel metal1 -574 553 -573 554 1 llama
<< end >>
