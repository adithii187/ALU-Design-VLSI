* SPICE3 file created from final_4.ext - technology: scmos

.option scale=0.09u

M1000 adsub_b2 a_n33840_n2871# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=347733 ps=33048
M1001 a_n29457_n8883# a_n30123_n8919# vdd w_n29547_n8685# pfet w=54 l=18
+  ad=2916 pd=216 as=635202 ps=50436
M1002 a_n28620_n5877# x2 vdd w_n28737_n5787# pfet w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1003 gnd comp_a1 a_n30123_n1953# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1004 AlessB a_n27072_n891# vdd w_n27144_n792# pfet w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1005 gnd D1 a_n30483_5634# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1006 D1 a_n35820_n12033# gnd Gnd nfet w=27 l=18
+  ad=13122 pd=1026 as=0 ps=0
M1007 a_n29565_6714# a_n29286_7263# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1008 a_n33840_n1935# D gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1009 a_n28620_n1548# x2 vdd w_n28737_n1458# pfet w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1010 AmoreB_2 a_n27954_n5094# vdd w_n27576_n5085# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1011 comp_a0 comp_b0 a_n30123_n3051# w_n29898_n3420# pfet w=63 l=18
+  ad=6318 pd=450 as=6804 ps=468
M1012 comp_b0 a_n30330_n12609# a_n30123_n12177# Gnd nfet w=54 l=18
+  ad=7290 pd=594 as=5832 ps=432
M1013 D1 a_n30690_9612# a_n30483_10044# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=8748 ps=648
M1014 a_n29637_6840# a_n29853_7128# vdd w_n29718_6822# pfet w=45 l=18
+  ad=3240 pd=234 as=0 ps=0
M1015 AmoreB_3 a_n28710_n4284# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1016 a_n30123_n1953# a_n30330_n2187# a_n30123_n1755# w_n29898_n2124# pfet w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1017 a_n29673_7749# adsub_a2 a_n29673_7947# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=8748 ps=648
M1018 a_n30483_3897# adsub_a0 a_n29673_3897# w_n29448_3528# pfet w=63 l=18
+  ad=10206 pd=702 as=10206 ps=702
M1019 a_n33822_n15822# D3 vdd w_n33912_n15849# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1020 gnd comp_a3 a_n30330_n9351# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1021 a_n30123_n6282# comp_a1 a_n30123_n6084# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1022 comp_a2 a_n33822_n8721# vdd w_n33444_n8712# pfet w=54 l=18
+  ad=6318 pd=450 as=0 ps=0
M1023 a_n30483_7749# a_n30690_7515# a_n30483_7947# w_n30258_7578# pfet w=63 l=18
+  ad=6804 pd=468 as=10206 ps=702
M1024 a_n28773_n7326# b0_not gnd Gnd nfet w=27 l=18
+  ad=2916 pd=270 as=0 ps=0
M1025 a_n31851_n13896# and_a3 vdd w_n31941_n13923# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1026 a_n29286_5148# carry0 a_n29286_5022# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1027 a0_not comp_a0 vdd w_n29268_n2817# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1028 adsub_b3 a_n33840_n2376# vdd w_n33462_n2367# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1029 a_n33822_n8226# a3 vdd w_n33912_n8253# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1030 a_n31851_n14373# and_b2 vdd w_n31941_n14400# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1031 a_n33822_n14508# D3 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1032 adsub_a1 a_n33840_n1278# vdd w_n33462_n1269# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1033 a_n30123_n4320# comp_a3 a_n30123_n4122# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1034 a_n33822_n10638# D2 vdd w_n33912_n10665# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1035 and_b2 a_n33822_n14877# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1036 a_n33840_n2871# b2 vdd w_n33930_n2898# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1037 a_n30123_n5265# a_n30330_n5499# a_n30123_n5067# w_n29898_n5436# pfet w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1038 a_n35685_n12600# s1 a_n35820_n12600# Gnd nfet w=27 l=18
+  ad=243 pd=72 as=3159 ps=288
M1039 a_n28323_n5166# a_n28782_n5094# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1040 a_n28791_7749# carry1 sum2 Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1041 a_n33822_n8847# D2 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1042 a_n28224_n6030# temp_more a_n28350_n6030# Gnd nfet w=27 l=18
+  ad=3159 pd=288 as=2916 ps=270
M1043 a_n33822_n12573# D3 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1044 gnd D1 a_n30483_3699# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1045 a_n33822_n15291# b1 vdd w_n33912_n15318# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1046 a_n28782_n765# a2_not vdd w_n28872_n792# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1047 vdd adsub_a2 a_n29880_7515# w_n29448_7578# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1048 gnd comp_a1 a_n30330_n6516# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1049 a_n29637_6723# a_n29853_7128# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1050 a_n30312_5085# adsub_a1 vdd w_n30402_5058# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1051 and_b1 a_n33822_n15291# vdd w_n33444_n15282# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1052 a3_not comp_a3 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1053 a_n30123_n7578# a_n30330_n7812# a_n30123_n7380# w_n29898_n7749# pfet w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1054 a_n27072_n5220# AmoreB_0 a_n26892_n5103# w_n27576_n5085# pfet w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1055 a_n29457_n9828# a_n30123_n9864# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1056 a_n28710_n4284# comp_a3 vdd w_n28800_n4311# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1057 a_n28152_n9981# a_n29457_n8883# gnd Gnd nfet w=27 l=18
+  ad=2916 pd=270 as=0 ps=0
M1058 a2_not comp_a2 vdd w_n29205_n675# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1059 x1 a_n30123_n6084# vdd w_n29547_n5850# pfet w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1060 a_n30123_n12375# comp_a0 a_n30123_n12177# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1061 a_n33822_n9135# D2 vdd w_n33912_n9162# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1062 a_n34407_n1233# D1 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1063 a_n35820_n12888# s0 a_n35703_n13014# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=729 ps=108
M1064 comp_b2 comp_a2 a_n30123_n9864# w_n29898_n10233# pfet w=63 l=18
+  ad=9720 pd=684 as=6804 ps=468
M1065 vdd comp_a2 a_n30330_n5499# w_n29898_n5436# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1066 D0 a_n35820_n11565# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1067 x1 a_n30123_n1755# vdd w_n29547_n1521# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1068 a_n35820_n12033# s1_not a_n35820_n12159# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1069 x3 a_n30123_n4122# vdd w_n29547_n3888# pfet w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1070 vdd comp_b2 a_n30330_n1170# w_n29898_n1107# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1071 a_n27756_n9981# a_n29457_n12141# a_n27882_n9981# Gnd nfet w=27 l=18
+  ad=3159 pd=288 as=2916 ps=270
M1072 a_n26892_n774# AlessB_1 a_n26982_n774# w_n27144_n792# pfet w=45 l=18
+  ad=3240 pd=234 as=3240 ps=234
M1073 a_n28791_9846# a_n28998_9612# sum3 w_n28566_9675# pfet w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1074 vdd a_n30285_n7686# a_n30330_n7812# w_n29898_n7749# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1075 comp_b0 comp_a0 a_n30123_n12177# w_n29898_n12546# pfet w=63 l=18
+  ad=9720 pd=684 as=6804 ps=468
M1076 comp_a0 a_n33822_n9666# gnd Gnd nfet w=27 l=18
+  ad=4374 pd=378 as=0 ps=0
M1077 vdd carry0 a_n28998_5400# w_n28566_5463# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1078 a_n30483_9846# a_n30690_9612# a_n30483_10044# w_n30258_9675# pfet w=63 l=18
+  ad=6804 pd=468 as=10206 ps=702
M1079 a_n33840_n864# D vdd w_n33930_n891# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1080 a_n33822_n11709# D2 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1081 a_n26811_n9945# k gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1082 vdd comp_b0 a_n30330_n3483# w_n29898_n3420# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1083 gnd comp_a0 a_n30330_n12609# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1084 a_n33822_n13887# a0 a_n33822_n14013# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1085 a_n28683_n891# comp_b2 a_n28782_n891# Gnd nfet w=27 l=9
+  ad=1215 pd=144 as=2430 ps=234
M1086 vdd D1 a_n28998_3465# w_n28566_3528# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1087 a_n33840_n3816# b0 a_n33840_n3942# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1088 a_n33822_n10143# b3 vdd w_n33912_n10170# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1089 gnd comp_a3 a_n30330_n4554# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1090 a_n30312_3150# adsub_a0 vdd w_n30402_3123# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1091 a_n28503_n2997# x2 a_n28647_n2997# Gnd nfet w=27 l=18
+  ad=2916 pd=270 as=3402 ps=306
M1092 comp_b3 a_n33822_n10143# vdd w_n33444_n10134# pfet w=54 l=18
+  ad=9720 pd=684 as=0 ps=0
M1093 a_n26892_n5103# AmoreB_1 a_n26982_n5103# w_n27576_n5085# pfet w=45 l=18
+  ad=0 pd=0 as=3240 ps=234
M1094 a_n31851_n13896# and_b3 vdd w_n31941_n13923# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1095 a_n30123_n9117# a_n30330_n9351# a_n30123_n8919# w_n29898_n9288# pfet w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1096 vdd a_n29673_10044# a_n28791_9846# w_n28566_9675# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1097 gnd adsub_a1 a_n29880_5400# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1098 a_n31851_n15237# and_a0 vdd w_n31941_n15264# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1099 a_n28377_n7326# x3 a_n28503_n7326# Gnd nfet w=27 l=18
+  ad=3159 pd=288 as=2916 ps=270
M1100 b0_not comp_b0 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1101 b1_not comp_b1 vdd w_n29214_n5850# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1102 a_n27072_n5220# AmoreB_3 gnd Gnd nfet w=27 l=18
+  ad=2916 pd=432 as=0 ps=0
M1103 a_n29637_8820# a_n29565_8811# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1104 a_n34407_n1233# D0 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1105 a_n33822_n12447# a3 vdd w_n33912_n12474# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1106 a_n28152_n9828# a_n29457_n9828# vdd w_n28260_n9846# pfet w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1107 a_n28773_n7173# b0_not vdd w_n28890_n7083# pfet w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1108 a_n28791_5634# a_n28998_5400# sum1 w_n28566_5463# pfet w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1109 and_oper_out2 a_n31851_n14373# vdd w_n31473_n14364# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1110 a0_not comp_a0 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1111 a_n33822_n14382# D3 vdd w_n33912_n14409# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1112 a1_not comp_a1 vdd w_n29214_n1521# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1113 gnd adsub_a0 a_n29880_3465# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1114 a_n30123_9# comp_b3 a_n30123_207# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1115 a_n33840_n369# a3 a_n33840_n495# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1116 a_n33840_n1809# a0 a_n33840_n1935# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1117 a_n33840_n2502# D gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1118 and_a3 a_n33822_n12447# vdd w_n33444_n12438# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1119 vdd adsub_b1 a_n30690_5400# w_n30258_5463# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1120 a_n33822_n11052# b1 a_n33822_n11178# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1121 gnd a_n30483_10044# a_n29673_9846# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1122 a_n27954_n765# x3 vdd w_n28044_n792# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1123 a_n29853_3078# a_n30312_3150# vdd w_n29934_3159# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1124 a_n30483_7947# adsub_a2 a_n29673_7947# w_n29448_7578# pfet w=63 l=18
+  ad=0 pd=0 as=10206 ps=702
M1125 vdd adsub_b0 a_n30690_3465# w_n30258_3528# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1126 a_n33822_n13068# D3 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1127 a_n29673_5634# adsub_a1 a_n29673_5832# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=8748 ps=648
M1128 a_n30312_3150# adsub_a0 a_n30312_3024# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1129 gnd carry0 a_n28998_5400# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1130 a_n28620_n5877# b1_not vdd w_n28737_n5787# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1131 vdd D1 a_n30483_9846# w_n30258_9675# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1132 a_n27954_n5094# x3 a_n27954_n5220# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1133 a_n30123_n12375# a_n30330_n12609# a_n30123_n12177# w_n29898_n12546# pfet w=63 l=18
+  ad=6804 pd=468 as=0 ps=0
M1134 a_n31851_n14022# and_a3 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1135 a_n28620_n1548# a1_not vdd w_n28737_n1458# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1136 b2_not comp_b2 vdd w_n29205_n5004# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1137 a_n28782_n765# comp_b2 vdd w_n28872_n792# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1138 a_n30483_5634# a_n30690_5400# a_n30483_5832# w_n30258_5463# pfet w=63 l=18
+  ad=6804 pd=468 as=10206 ps=702
M1139 x1 a_n30123_n6084# gnd Gnd nfet w=27 l=18
+  ad=2916 pd=324 as=0 ps=0
M1140 gnd D1 a_n28998_3465# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1141 gnd adsub_b3 a_n30690_9612# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1142 comp_b2 a_n30330_n5499# a_n30123_n5067# Gnd nfet w=54 l=18
+  ad=7290 pd=594 as=5832 ps=432
M1143 gnd a_n29673_10044# a_n28791_9846# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1144 a_n29286_5148# carry0 vdd w_n29376_5121# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1145 vdd comp_b3 a_n30123_n9117# w_n29898_n9288# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1146 adsub_a0 a_n33840_n1809# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1147 k a_n28152_n9828# gnd Gnd nfet w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
M1148 a_n33822_n8721# a2 a_n33822_n8847# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1149 a_n28791_3699# a_n28998_3465# sum0 w_n28566_3528# pfet w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1150 a_n28620_n5877# x3 a_n28224_n6030# Gnd nfet w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1151 a_n29286_5022# a_n29673_5832# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1152 a_n29853_3078# a_n30312_3150# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1153 a_n35820_n12888# s1 vdd w_n35910_n12915# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1154 a_n33822_n8721# D2 vdd w_n33912_n8748# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1155 x3 a_n30123_n4122# gnd Gnd nfet w=27 l=18
+  ad=2916 pd=324 as=0 ps=0
M1156 a_n28791_5634# carry0 sum1 Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1157 a_n29673_5832# carry0 sum1 w_n28566_5463# pfet w=63 l=18
+  ad=10206 pd=702 as=0 ps=0
M1158 vdd comp_a0 a_n30330_n12609# w_n29898_n12546# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1159 carry1 a_n29637_4608# vdd w_n29718_4707# pfet w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1160 a_n27018_n5103# AmoreB_3 a_n27072_n5103# w_n27576_n5085# pfet w=45 l=18
+  ad=810 pd=126 as=1620 ps=162
M1161 and_oper_out1 a_n31851_n14769# vdd w_n31473_n14760# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1162 comp_a0 a_n30330_n3483# a_n30123_n3051# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1163 a_n33822_n11583# D2 vdd w_n33912_n11610# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1164 adsub_b1 a_n33840_n3285# vdd w_n33462_n3276# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1165 and_b0 a_n33822_n15822# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1166 a_n33822_n9135# a1 vdd w_n33912_n9162# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1167 a_n30483_10044# a_n29880_9612# a_n29673_10044# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=8748 ps=648
M1168 a_n31851_n14769# and_a1 vdd w_n31941_n14796# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1169 a_n33822_n15417# D3 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1170 a_n30123_n11079# comp_a1 a_n30123_n10881# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1171 a_n29673_3699# adsub_a0 a_n29673_3897# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=8748 ps=648
M1172 a_n30123_n1953# comp_b1 a_n30123_n1755# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1173 a_n30312_5085# a_n30483_5832# vdd w_n30402_5058# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1174 carry0 a_n29637_2673# vdd w_n29718_2772# pfet w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1175 a_n31851_n15237# and_b0 vdd w_n31941_n15264# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1176 a_n33822_n9792# D2 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1177 a_n28494_n6030# comp_a1 a_n28620_n6030# Gnd nfet w=27 l=18
+  ad=3402 pd=306 as=2916 ps=270
M1178 comp_a3 a_n33822_n8226# gnd Gnd nfet w=27 l=18
+  ad=4374 pd=378 as=0 ps=0
M1179 AlessB_0 a_n28773_n2844# gnd Gnd nfet w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
M1180 and_oper_out3 a_n31851_n13896# vdd w_n31473_n13887# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1181 gnd comp_b3 a_n30330_n225# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1182 a_n33822_n13482# D3 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1183 a_n30483_5832# a_n29880_5400# a_n29673_5832# Gnd nfet w=54 l=18
+  ad=8748 pd=648 as=0 ps=0
M1184 a_n33822_n13887# D3 vdd w_n33912_n13914# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1185 a_n33822_n10269# D2 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1186 a_n30483_3699# a_n30690_3465# a_n30483_3897# w_n30258_3528# pfet w=63 l=18
+  ad=6804 pd=468 as=0 ps=0
M1187 a_n28152_n9828# temp a_n27756_n9981# Gnd nfet w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1188 a_n28773_n7173# x3 vdd w_n28890_n7083# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1189 a_n35820_n12033# s1_not vdd w_n35910_n12060# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1190 b1_not comp_b1 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1191 gnd D1 a_n30483_7749# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1192 a_n35820_n11691# s0_not gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1193 D1 adsub_b1 a_n30483_5832# w_n30258_5463# pfet w=63 l=18
+  ad=16524 pd=1152 as=0 ps=0
M1194 a_n29286_3213# D1 vdd w_n29376_3186# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1195 a_n28224_n1701# temp_less a_n28350_n1701# Gnd nfet w=27 l=18
+  ad=3159 pd=288 as=2916 ps=270
M1196 a_n29286_3213# D1 a_n29286_3087# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1197 a_n26811_n9819# equals_d a_n26811_n9945# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1198 carry1 a_n29637_4608# gnd Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1199 a_n30123_n5265# comp_a2 a_n30123_n5067# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1200 a_n28791_3699# D1 sum0 Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1201 a_n29637_8820# a_n29853_9225# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1202 a_n29673_3897# D1 sum0 w_n28566_3528# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1203 D2 a_n35820_n12474# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1204 AlessB_2 a_n27954_n765# vdd w_n27576_n756# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1205 adsub_a3 a_n33840_n369# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1206 carry0 a_n29637_2673# gnd Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1207 adsub_a2 a_n33840_n864# vdd w_n33462_n855# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1208 a_n29673_5832# a_n28998_5400# sum1 Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1209 vdd comp_b1 a_n30123_n6282# w_n29898_n6453# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1210 a_n31851_n13896# and_b3 a_n31851_n14022# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1211 a_n30123_n7578# a_n30285_n7686# a_n30123_n7380# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1212 a_n33822_n10638# b2 a_n33822_n10764# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1213 a_n28773_n2844# x2 vdd w_n28890_n2754# pfet w=54 l=18
+  ad=17496 pd=1188 as=0 ps=0
M1214 a_n28773_n7173# a_n30285_n7686# a_n28377_n7326# Gnd nfet w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1215 a_n27954_n5094# x3 vdd w_n28044_n5121# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1216 vdd a_n30483_5832# a_n29673_5634# w_n29448_5463# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1217 a_n26982_n5103# AmoreB_3 a_n27018_n5103# w_n27576_n5085# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1218 a_n30312_3150# a_n30483_3897# vdd w_n30402_3123# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1219 gnd comp_b1 a_n30123_n11079# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1220 a_n29673_10044# a_n28998_9612# sum3 Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1221 comp_a2 a_n30330_n1170# a_n30123_n738# Gnd nfet w=54 l=18
+  ad=4374 pd=378 as=5832 ps=432
M1222 a_n33840_n2376# b3 a_n33840_n2502# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1223 comp_b2 a_n33822_n10638# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1224 a_n28323_n837# a_n28782_n765# vdd w_n28404_n756# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1225 a_n30483_3897# a_n29880_3465# a_n29673_3897# Gnd nfet w=54 l=18
+  ad=8748 pd=648 as=0 ps=0
M1226 a_n29457_n12141# a_n30123_n12177# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1227 comp_b2 a_n30330_n10296# a_n30123_n9864# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1228 AmoreB_1 a_n28620_n5877# vdd w_n28737_n5787# pfet w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1229 gnd comp_a2 a_n30330_n5499# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1230 vdd comp_b3 a_n30123_n4320# w_n29898_n4491# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1231 a_n29637_8820# a_n29565_8811# a_n29637_8937# w_n29718_8919# pfet w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1232 a_n33822_n11052# b1 vdd w_n33912_n11079# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1233 gnd comp_a2 a_n30330_n10296# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1234 AlessB_1 a_n28620_n1548# vdd w_n28737_n1458# pfet w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1235 gnd comp_b2 a_n30330_n1170# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1236 comp_a2 comp_b2 a_n30123_n738# w_n29898_n1107# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1237 AequalsB a_n26811_n9819# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1238 a_n28647_n7326# x1 a_n28773_n7326# Gnd nfet w=27 l=18
+  ad=3402 pd=306 as=0 ps=0
M1239 comp_b1 a_n33822_n11052# vdd w_n33444_n11043# pfet w=54 l=18
+  ad=9720 pd=684 as=0 ps=0
M1240 a_n30483_7749# adsub_b2 a_n30483_7947# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=8748 ps=648
M1241 vdd carry1 a_n28998_7515# w_n28566_7578# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1242 a_n30312_7200# adsub_a2 vdd w_n30402_7173# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1243 a_n33840_n495# D gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1244 D1 adsub_b0 a_n30483_3897# w_n30258_3528# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1245 a_n30312_7200# adsub_a2 a_n30312_7074# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1246 gnd a_n30285_n7686# a_n30330_n7812# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1247 x2 a_n30123_n5067# vdd w_n29547_n4833# pfet w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1248 a_n30123_9# a_n30330_n225# a_n30123_207# w_n29898_n162# pfet w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1249 AlessB_3 a_n28710_45# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1250 a_n31851_n14769# and_b1 vdd w_n31941_n14796# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1251 a_n30123_n11079# a_n30330_n11313# a_n30123_n10881# w_n29898_n11250# pfet w=63 l=18
+  ad=6804 pd=468 as=6804 ps=468
M1252 a_n27954_n891# a_n28323_n837# gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1253 a_n33822_n13356# a1 vdd w_n33912_n13383# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1254 a_n29673_9846# a_n29880_9612# a_n29673_10044# w_n29448_9675# pfet w=63 l=18
+  ad=6804 pd=468 as=10206 ps=702
M1255 gnd comp_a2 a_n30123_n936# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1256 gnd comp_b0 a_n30330_n3483# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1257 a_n27018_n774# AlessB_3 a_n27072_n774# w_n27144_n792# pfet w=45 l=18
+  ad=810 pd=126 as=1620 ps=162
M1258 a_n33822_n15291# D3 vdd w_n33912_n15318# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1259 a_n33840_n3411# D gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1260 and_a1 a_n33822_n13356# vdd w_n33444_n13347# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1261 a_n33840_n3816# D vdd w_n33930_n3843# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1262 a_n30312_3024# a_n30483_3897# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1263 a_n35820_n11565# s1_not vdd w_n35910_n11592# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1264 a_n29673_3897# a_n28998_3465# sum0 Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1265 x2 a_n30123_n738# gnd Gnd nfet w=27 l=18
+  ad=2916 pd=324 as=0 ps=0
M1266 and_oper_out0 a_n31851_n15237# vdd w_n31473_n15228# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1267 gnd adsub_a2 a_n29880_7515# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1268 vdd a_n30483_3897# a_n29673_3699# w_n29448_3528# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1269 AlessB_3 a_n28710_45# vdd w_n28332_54# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1270 a_n28710_45# comp_b3 a_n28611_n81# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=1215 ps=144
M1271 vdd comp_a2 a_n30123_n936# w_n29898_n1107# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1272 a_n30123_n9117# comp_a3 a_n30123_n8919# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=5832 ps=432
M1273 adsub_b2 a_n33840_n2871# vdd w_n33462_n2862# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1274 a_n28350_n6030# x2 a_n28494_n6030# Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1275 x0 a_n30123_n3051# vdd w_n29547_n2817# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1276 a_n33822_n8721# a2 vdd w_n33912_n8748# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1277 a_n29853_7128# a_n30312_7200# vdd w_n29934_7209# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1278 D1 a_n35820_n12033# vdd w_n35442_n12024# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1279 a_n35820_n13014# s1 gnd Gnd nfet w=27 l=18
+  ad=2673 pd=252 as=0 ps=0
M1280 vdd adsub_b2 a_n30690_7515# w_n30258_7578# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1281 a_n33840_n1404# D gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1282 D a_n34407_n1233# gnd Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1283 a_n33840_n1809# D vdd w_n33930_n1836# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1284 a_n29286_5148# a_n29673_5832# vdd w_n29376_5121# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1285 a_n28611_n4410# comp_a3 a_n28710_n4410# Gnd nfet w=27 l=9
+  ad=1215 pd=144 as=2430 ps=234
M1286 a_n35820_n12159# s0 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1287 AmoreB_3 a_n28710_n4284# vdd w_n28332_n4275# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1288 a_n35820_n12474# s1 a_n35685_n12600# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1289 a_n29565_8811# a_n29286_9360# vdd w_n28908_9369# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1290 a_n33822_n9666# a0 a_n33822_n9792# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1291 gnd carry1 a_n28998_7515# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1292 adsub_b0 a_n33840_n3816# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1293 s0_not s0 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1294 vdd comp_b1 a_n30123_n11079# w_n29898_n11250# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1295 a_n27882_n9981# a_n29457_n10845# a_n28026_n9981# Gnd nfet w=27 l=18
+  ad=0 pd=0 as=3402 ps=306
M1296 a_n33822_n14013# D3 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1297 a_n33822_n14877# b2 vdd w_n33912_n14904# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1298 AlessB_0 a_n28773_n2844# vdd w_n28890_n2754# pfet w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1299 a_n28773_n7173# a_n30285_n7686# vdd w_n28890_n7083# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1300 a_n33822_n10143# D2 vdd w_n33912_n10170# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1301 a_n29853_7128# a_n30312_7200# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1302 and_b3 a_n33822_n14382# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1303 a3_not comp_a3 vdd w_n29178_135# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1304 and_b2 a_n33822_n14877# vdd w_n33444_n14868# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1305 a_n30483_9846# adsub_b3 a_n30483_10044# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1306 a_n28773_n2997# a0_not gnd Gnd nfet w=27 l=18
+  ad=2916 pd=270 as=0 ps=0
M1307 a_n29286_7263# carry1 vdd w_n29376_7236# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1308 vdd comp_a2 a_n30330_n10296# w_n29898_n10233# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1309 a_n33822_n8352# D2 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1310 a_n28323_n5166# a_n28782_n5094# vdd w_n28404_n5085# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1311 a_n28620_n1548# x3 a_n28224_n1701# Gnd nfet w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1312 s1_not s1 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1313 vdd comp_b3 a_n30330_n225# w_n29898_n162# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1314 gnd comp_b3 a_n30123_n9117# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1315 a_n33822_n12447# D3 vdd w_n33912_n12474# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1316 a_n29565_8811# a_n29286_9360# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1317 a_n29673_7947# carry1 sum2 w_n28566_7578# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1318 carry2 a_n29637_6723# vdd w_n29718_6822# pfet w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1319 a_n29286_3213# a_n29673_3897# vdd w_n29376_3186# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1320 a_n28773_n7173# x1 vdd w_n28890_n7083# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1321 a_n27954_n5220# a_n28323_n5166# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1322 a_n29457_n9828# a_n30123_n9864# vdd w_n29547_n9630# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1323 a_n29286_3087# a_n29673_3897# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1324 a_n33822_n11178# D2 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1325 x2 a_n30123_n5067# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1326 a_n29637_8937# a_n29853_9225# vdd w_n29718_8919# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1327 gnd adsub_b1 a_n30690_5400# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1328 a_n28152_n9828# a_n29457_n8883# vdd w_n28260_n9846# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1329 a_n34407_n1233# D1 a_n34407_n1116# w_n34488_n1134# pfet w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1330 comp_b2 a_n33822_n10638# vdd w_n33444_n10629# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1331 a_n30123_n3249# a_n30330_n3483# a_n30123_n3051# w_n29898_n3420# pfet w=63 l=18
+  ad=6804 pd=468 as=0 ps=0
M1332 a_n28494_n1701# comp_b1 a_n28620_n1701# Gnd nfet w=27 l=18
+  ad=3402 pd=306 as=2916 ps=270
M1333 D0 a_n35820_n11565# vdd w_n35442_n11556# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1334 a_n29457_n10845# a_n30123_n10881# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1335 b3_not comp_b3 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1336 a_n29457_n7344# a_n30123_n7380# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1337 gnd adsub_b0 a_n30690_3465# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1338 a_n27072_n891# AlessB_3 gnd Gnd nfet w=27 l=18
+  ad=2916 pd=432 as=0 ps=0
M1339 a_n30483_7947# a_n29880_7515# a_n29673_7947# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1340 a_n33822_n12942# a2 vdd w_n33912_n12969# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1341 a_n29286_7263# carry1 a_n29286_7137# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1342 x0 a_n30123_n3051# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1343 and_a2 a_n33822_n12942# vdd w_n33444_n12933# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1344 gnd D1 a_n30483_9846# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1345 a_n28152_n9828# a_n29457_n12141# vdd w_n28260_n9846# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1346 comp_b0 a_n30285_n7686# a_n30123_n7380# w_n29898_n7749# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1347 comp_a0 a_n33822_n9666# vdd w_n33444_n9657# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1348 a_n33822_n15822# b0 a_n33822_n15948# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1349 comp_a1 a_n33822_n9135# gnd Gnd nfet w=27 l=18
+  ad=4374 pd=378 as=0 ps=0
M1350 D1 adsub_b2 a_n30483_7947# w_n30258_7578# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1351 a_n33840_n2376# D vdd w_n33930_n2403# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1352 carry2 a_n29637_6723# gnd Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1353 a_n30483_5634# adsub_b1 a_n30483_5832# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1354 comp_b0 a_n33822_n11583# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1355 a_n26811_n9819# k vdd w_n26901_n9846# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1356 vdd adsub_a3 a_n29880_9612# w_n29448_9675# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1357 a_n33840_n3285# b1 a_n33840_n3411# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1358 a_n27072_n891# AlessB_0 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1359 a_n33840_n3816# b0 vdd w_n33930_n3843# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1360 a_n30312_7200# a_n30483_7947# vdd w_n30402_7173# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1361 a_n27072_n891# AlessB_2 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1362 a_n30312_7074# a_n30483_7947# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1363 a_n29673_7947# a_n28998_7515# sum2 Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1364 b0_not comp_b0 vdd w_n29268_n7146# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1365 and_a0 a_n33822_n13887# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1366 gnd comp_b1 a_n30123_n6282# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1367 a_n34407_n1116# D0 vdd w_n34488_n1134# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1368 a_n28683_n5220# comp_a2 a_n28782_n5220# Gnd nfet w=27 l=9
+  ad=1215 pd=144 as=2430 ps=234
M1369 a_n33840_n1278# a1 a_n33840_n1404# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1370 a_n28377_n2997# x3 a_n28503_n2997# Gnd nfet w=27 l=18
+  ad=3159 pd=288 as=0 ps=0
M1371 a_n33840_n369# a3 vdd w_n33930_n396# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1372 a_n33840_n1809# a0 vdd w_n33930_n1836# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1373 vdd comp_a0 a_n30123_n3249# w_n29898_n3420# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1374 AlessB a_n27072_n891# gnd Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1375 a_n29457_n8883# a_n30123_n8919# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1376 gnd comp_b3 a_n30123_n4320# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1377 x3 a_n30123_207# vdd w_n29547_441# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1378 vdd comp_b1 a_n30330_n2187# w_n29898_n2124# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1379 a_n30312_5085# adsub_a1 a_n30312_4959# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1380 a_n28710_n81# a3_not gnd Gnd nfet w=27 l=18
+  ad=2430 pd=234 as=0 ps=0
M1381 a_n35820_n12033# s0 vdd w_n35910_n12060# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1382 a_n35820_n12474# s1 vdd w_n35910_n12501# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1383 AmoreB_2 a_n27954_n5094# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1384 vdd comp_b2 a_n30123_n5265# w_n29898_n5436# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1385 comp_b3 comp_a3 a_n30123_n8919# w_n29898_n9288# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1386 a_n28620_n6030# b1_not gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1387 a_n30483_3699# adsub_b0 a_n30483_3897# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1388 a_n30312_9297# adsub_a3 a_n30312_9171# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1389 a_n28782_n5220# b2_not gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1390 a_n27954_n5094# a_n28323_n5166# vdd w_n28044_n5121# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1391 vdd a_n30483_7947# a_n29673_7749# w_n29448_7578# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1392 vdd comp_b0 a_n30123_n7578# w_n29898_n7749# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1393 D1 a_n30690_5400# a_n30483_5832# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1394 vdd a_n29673_5832# a_n28791_5634# w_n28566_5463# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1395 a_n33822_n14877# b2 a_n33822_n15003# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1396 a_n29637_4608# a_n29565_4599# a_n29637_4725# w_n29718_4707# pfet w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1397 comp_a2 a_n33822_n8721# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1398 a_n28611_n81# comp_b3 a_n28710_n81# Gnd nfet w=27 l=9
+  ad=0 pd=0 as=0 ps=0
M1399 a_n33822_n8226# a3 a_n33822_n8352# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1400 gnd comp_b0 a_n30123_n12375# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1401 adsub_b3 a_n33840_n2376# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1402 D3 a_n35820_n12888# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1403 a_n28350_n1701# x2 a_n28494_n1701# Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1404 adsub_a0 a_n33840_n1809# vdd w_n33462_n1800# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1405 a_n33822_n10764# D2 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1406 x3 a_n30123_207# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1407 a_n28773_n2844# a0_not vdd w_n28890_n2754# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1408 a_n29637_2673# a_n29565_2664# a_n29637_2790# w_n29718_2772# pfet w=45 l=18
+  ad=1215 pd=144 as=3240 ps=234
M1409 a_n29853_9225# a_n30312_9297# vdd w_n29934_9306# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1410 k a_n28152_n9828# vdd w_n28260_n9846# pfet w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1411 a_n30123_n10062# a_n30330_n10296# a_n30123_n9864# w_n29898_n10233# pfet w=63 l=18
+  ad=6804 pd=468 as=0 ps=0
M1412 a_n28782_n891# a2_not gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1413 gnd a_n30483_5832# a_n29673_5634# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1414 and_a2 a_n33822_n12942# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1415 a_n27072_n5220# AmoreB_2 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1416 a_n28620_n5877# temp_more vdd w_n28737_n5787# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1417 a_n29286_7263# a_n29673_7947# vdd w_n29376_7236# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1418 a_n29673_10044# carry2 sum3 w_n28566_9675# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1419 a_n28782_n5094# comp_a2 a_n28683_n5220# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1420 and_b0 a_n33822_n15822# vdd w_n33444_n15813# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1421 a_n33822_n11052# D2 vdd w_n33912_n11079# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1422 and_b1 a_n33822_n15291# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1423 a_n28620_n1548# temp_less vdd w_n28737_n1458# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1424 vdd D1 a_n30483_5634# w_n30258_5463# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1425 a2_not comp_a2 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1426 D1 adsub_b3 a_n30483_10044# w_n30258_9675# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1427 vdd comp_a3 a_n30123_9# w_n29898_n162# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1428 comp_a3 a_n33822_n8226# vdd w_n33444_n8217# pfet w=54 l=18
+  ad=6318 pd=450 as=0 ps=0
M1429 a_n33822_n9261# D2 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1430 a_n29637_4608# a_n29565_4599# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1431 a_n33822_n9666# D2 vdd w_n33912_n9693# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1432 AmoreB a_n27072_n5220# gnd Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1433 D1 a_n30690_3465# a_n30483_3897# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1434 a_n33822_n13356# D3 vdd w_n33912_n13383# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1435 vdd a_n29673_3897# a_n28791_3699# w_n28566_3528# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1436 a_n29673_7749# a_n29880_7515# a_n29673_7947# w_n29448_7578# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1437 x1 a_n30123_n1755# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1438 gnd a_n29673_5832# a_n28791_5634# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1439 a_n29637_2673# a_n29565_2664# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=216 as=0 ps=0
M1440 comp_b1 comp_a1 a_n30123_n6084# w_n29898_n6453# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1441 a_n29853_9225# a_n30312_9297# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1442 a_n33840_n2376# b3 vdd w_n33930_n2403# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1443 a_n28152_n9828# temp vdd w_n28260_n9846# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1444 a_n35820_n11565# s0_not vdd w_n35910_n11592# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1445 a_n27072_n891# AlessB_1 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1446 a_n33822_n15822# b0 vdd w_n33912_n15849# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1447 a_n29286_9360# carry2 vdd w_n29376_9333# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1448 a_n29565_4599# a_n29286_5148# vdd w_n28908_5157# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1449 comp_b1 a_n30330_n11313# a_n30123_n10881# Gnd nfet w=54 l=18
+  ad=7290 pd=594 as=0 ps=0
M1450 comp_a1 comp_b1 a_n30123_n1755# w_n29898_n2124# pfet w=63 l=18
+  ad=6318 pd=450 as=0 ps=0
M1451 a_n29673_9846# adsub_a3 a_n29673_10044# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1452 a_n29286_7137# a_n29673_7947# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1453 a_n26811_n9819# equals_d vdd w_n26901_n9846# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1454 a_n33840_n2997# D gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1455 a_n28503_n7326# x2 a_n28647_n7326# Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1456 gnd a_n30483_3897# a_n29673_3699# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1457 comp_a3 a_n30330_n225# a_n30123_207# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1458 comp_b3 comp_a3 a_n30123_n4122# w_n29898_n4491# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1459 D2 a_n35820_n12474# vdd w_n35442_n12465# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1460 adsub_a3 a_n33840_n369# vdd w_n33462_n360# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1461 a_n33822_n14382# b3 a_n33822_n14508# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1462 a_n28782_n5094# b2_not vdd w_n28872_n5121# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1463 gnd adsub_b2 a_n30690_7515# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1464 a_n33822_n10638# b2 vdd w_n33912_n10665# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1465 vdd D1 a_n30483_3699# w_n30258_3528# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1466 comp_b3 a_n33822_n10143# gnd Gnd nfet w=27 l=18
+  ad=7290 pd=594 as=0 ps=0
M1467 a_n35820_n12600# s0_not gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1468 a_n31851_n15363# and_a0 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1469 a_n33840_n3285# D vdd w_n33930_n3312# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1470 a_n28026_n9981# a_n29457_n9828# a_n28152_n9981# Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1471 vdd comp_b0 a_n30123_n12375# w_n29898_n12546# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1472 a_n33822_n12447# a3 a_n33822_n12573# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1473 vdd comp_a1 a_n30123_n1953# w_n29898_n2124# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1474 a_n28710_45# a3_not vdd w_n28800_18# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1475 AmoreB_1 a_n28620_n5877# gnd Gnd nfet w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
M1476 a_n30123_n3249# comp_b0 a_n30123_n3051# Gnd nfet w=54 l=18
+  ad=5832 pd=432 as=0 ps=0
M1477 a_n29457_n12141# a_n30123_n12177# vdd w_n29547_n11943# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1478 a_n28773_n2844# comp_b0 a_n28377_n2997# Gnd nfet w=27 l=18
+  ad=3645 pd=324 as=0 ps=0
M1479 a_n28773_n2844# x3 vdd w_n28890_n2754# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1480 a_n29565_4599# a_n29286_5148# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1481 and_oper_out2 a_n31851_n14373# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1482 a_n31851_n14499# and_a2 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1483 a1_not comp_a1 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1484 a_n29286_9360# carry2 a_n29286_9234# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1485 and_a3 a_n33822_n12447# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1486 gnd a_n29673_3897# a_n28791_3699# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1487 a_n33822_n14877# D3 vdd w_n33912_n14904# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1488 AequalsB a_n26811_n9819# vdd w_n26433_n9810# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1489 a_n33840_n864# a2 a_n33840_n990# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=3888 ps=342
M1490 a_n27954_n765# x3 a_n27954_n891# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1491 a_n33840_n369# D vdd w_n33930_n396# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1492 a_n33840_n1278# D vdd w_n33930_n1305# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1493 vdd comp_a3 a_n30330_n9351# w_n29898_n9288# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1494 comp_b0 a_n30330_n7812# a_n30123_n7380# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1495 a_n29637_4725# a_n29853_5013# vdd w_n29718_4707# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1496 a_n29565_2664# a_n29286_3213# vdd w_n28908_3222# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1497 a_n30123_n6282# a_n30330_n6516# a_n30123_n6084# w_n29898_n6453# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1498 carry3 a_n29637_8820# gnd Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1499 a_n27954_n765# a_n28323_n837# vdd w_n28044_n792# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1500 a_n30312_4959# a_n30483_5832# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1501 a_n28782_n5094# comp_a2 vdd w_n28872_n5121# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1502 a_n28647_n2997# x1 a_n28773_n2997# Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1503 a_n28791_9846# carry2 sum3 Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1504 a_n28710_n4410# b3_not gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1505 a_n30312_9297# adsub_a3 vdd w_n30402_9270# pfet w=45 l=18
+  ad=4455 pd=378 as=0 ps=0
M1506 a_n29637_2790# a_n29853_3078# vdd w_n29718_2772# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1507 x2 a_n30123_n738# vdd w_n29547_n504# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1508 a_n30312_9171# a_n30483_10044# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1509 a_n28782_n765# comp_b2 a_n28683_n891# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1510 D3 a_n35820_n12888# vdd w_n35442_n12879# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1511 a_n30123_n4320# a_n30330_n4554# a_n30123_n4122# w_n29898_n4491# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1512 b2_not comp_b2 gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1513 a_n33822_n11583# b0 a_n33822_n11709# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1514 vdd comp_a1 a_n30330_n6516# w_n29898_n6453# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1515 comp_b1 comp_a1 a_n30123_n10881# w_n29898_n11250# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1516 gnd comp_a3 a_n30123_9# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1517 a_n28620_n5877# x3 vdd w_n28737_n5787# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1518 a_n27072_n5103# AmoreB_2 vdd w_n27576_n5085# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1519 a_n29565_2664# a_n29286_3213# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1520 D a_n34407_n1233# vdd w_n34488_n1134# pfet w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1521 vdd adsub_a1 a_n29880_5400# w_n29448_5463# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1522 gnd comp_a0 a_n30123_n3249# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1523 a_n29637_4608# a_n29853_5013# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1524 a_n33822_n12942# D3 vdd w_n33912_n12969# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1525 a_n30123_n936# comp_b2 a_n30123_n738# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1526 gnd comp_a1 a_n30330_n11313# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1527 a_n28620_n1548# x3 vdd w_n28737_n1458# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1528 gnd comp_b1 a_n30330_n2187# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1529 a_n28620_n1701# a1_not gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1530 vdd carry2 a_n28998_9612# w_n28566_9675# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1531 AmoreB_0 a_n28773_n7173# gnd Gnd nfet w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
M1532 vdd adsub_a0 a_n29880_3465# w_n29448_3528# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1533 and_oper_out1 a_n31851_n14769# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1534 a_n31851_n14895# and_a1 gnd Gnd nfet w=27 l=18
+  ad=3888 pd=342 as=0 ps=0
M1535 a_n28773_n7173# x2 vdd w_n28890_n7083# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1536 a_n33822_n9135# a1 a_n33822_n9261# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1537 gnd comp_b2 a_n30123_n5265# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1538 adsub_b0 a_n33840_n3816# vdd w_n33462_n3807# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1539 a_n33822_n9666# a0 vdd w_n33912_n9693# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1540 a_n29637_2673# a_n29853_3078# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1541 adsub_b1 a_n33840_n3285# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1542 a_n33822_n15948# D3 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1543 comp_b3 a_n30330_n9351# a_n30123_n8919# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1544 s0_not s0 vdd w_n36243_n12096# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1545 gnd comp_b2 a_n30123_n10062# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=5832 ps=432
M1546 AmoreB a_n27072_n5220# vdd w_n27576_n5085# pfet w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1547 a_n33822_n14382# b3 vdd w_n33912_n14409# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1548 a_n31851_n15237# and_b0 a_n31851_n15363# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1549 a_n30123_n936# a_n30330_n1170# a_n30123_n738# w_n29898_n1107# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1550 vdd a_n30483_10044# a_n29673_9846# w_n29448_9675# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1551 D1 a_n30690_7515# a_n30483_7947# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1552 a_n28620_n5877# comp_a1 vdd w_n28737_n5787# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1553 a_n35703_n13014# s0 a_n35820_n13014# Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1554 and_b3 a_n33822_n14382# vdd w_n33444_n14373# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1555 a_n29637_6723# a_n29565_6714# a_n29637_6840# w_n29718_6822# pfet w=45 l=18
+  ad=1215 pd=144 as=0 ps=0
M1556 and_oper_out3 a_n31851_n13896# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1557 gnd comp_b0 a_n30123_n7578# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1558 a_n28152_n9828# a_n29457_n10845# vdd w_n28260_n9846# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1559 a_n29673_5634# a_n29880_5400# a_n29673_5832# w_n29448_5463# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1560 a_n28620_n1548# comp_b1 vdd w_n28737_n1458# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1561 gnd adsub_a3 a_n29880_9612# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1562 a_n31851_n14373# and_b2 a_n31851_n14499# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1563 a_n33822_n8226# D2 vdd w_n33912_n8253# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1564 adsub_a1 a_n33840_n1278# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1565 a_n33822_n12942# a2 a_n33822_n13068# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1566 s1_not s1 vdd w_n36234_n12420# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1567 a_n33840_n2871# b2 a_n33840_n2997# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1568 a_n33840_n2871# D vdd w_n33930_n2898# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1569 a_n30123_n10062# comp_a2 a_n30123_n9864# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1570 vdd adsub_b3 a_n30690_9612# w_n30258_9675# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1571 vdd comp_a3 a_n30330_n4554# w_n29898_n4491# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1572 a_n29286_9360# a_n29673_10044# vdd w_n29376_9333# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1573 AlessB_2 a_n27954_n765# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1574 a_n27072_n5220# AmoreB_0 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1575 vdd a_n29673_7947# a_n28791_7749# w_n28566_7578# pfet w=63 l=18
+  ad=0 pd=0 as=6804 ps=468
M1576 adsub_a2 a_n33840_n864# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1577 a_n33840_n3285# b1 vdd w_n33930_n3312# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1578 a_n28710_n4284# b3_not vdd w_n28800_n4311# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1579 a_n35820_n12474# s0_not vdd w_n35910_n12501# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1580 gnd carry2 a_n28998_9612# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=2916 ps=216
M1581 a_n29637_6723# a_n29565_6714# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1582 comp_a3 comp_b3 a_n30123_207# w_n29898_n162# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1583 b3_not comp_b3 vdd w_n29178_n4194# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1584 a_n29457_n10845# a_n30123_n10881# vdd w_n29547_n10647# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1585 a_n35820_n12888# s0 vdd w_n35910_n12915# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1586 a_n29457_n7344# a_n30123_n7380# vdd w_n29547_n7146# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1587 a_n30483_10044# adsub_a3 a_n29673_10044# w_n29448_9675# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1588 a_n29853_5013# a_n30312_5085# vdd w_n29934_5094# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1589 a_n26982_n774# AlessB_3 a_n27018_n774# w_n27144_n792# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1590 a_n28773_n2844# comp_b0 vdd w_n28890_n2754# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1591 a_n31851_n14373# and_a2 vdd w_n31941_n14400# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1592 a_n28323_n837# a_n28782_n765# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1593 a_n33822_n15003# D3 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1594 a_n29673_3699# a_n29880_3465# a_n29673_3897# w_n29448_3528# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1595 a_n33840_n864# a2 vdd w_n33930_n891# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1596 a_n33822_n11583# b0 vdd w_n33912_n11610# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1597 comp_a1 a_n33822_n9135# vdd w_n33444_n9126# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1598 gnd a_n30483_7947# a_n29673_7749# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1599 comp_b1 a_n30330_n6516# a_n30123_n6084# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1600 a_n33840_n1278# a1 vdd w_n33930_n1305# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1601 a_n33822_n15291# b1 a_n33822_n15417# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1602 a_n29565_6714# a_n29286_7263# vdd w_n28908_7272# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1603 vdd comp_a1 a_n30330_n11313# w_n29898_n11250# pfet w=63 l=18
+  ad=0 pd=0 as=3402 ps=234
M1604 comp_b0 a_n33822_n11583# vdd w_n33444_n11574# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1605 a_n30483_5832# adsub_a1 a_n29673_5832# w_n29448_5463# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1606 comp_b1 a_n33822_n11052# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1607 a_n29286_9234# a_n29673_10044# gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1608 comp_a1 a_n30330_n2187# a_n30123_n1755# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1609 a_n33840_n990# D gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1610 a_n31851_n14769# and_b1 a_n31851_n14895# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1611 a_n28710_n4284# comp_a3 a_n28611_n4410# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1612 vdd D1 a_n30483_7749# w_n30258_7578# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1613 a_n33822_n13356# a1 a_n33822_n13482# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1614 a_n27072_n891# AlessB_0 a_n26892_n774# w_n27144_n792# pfet w=45 l=18
+  ad=1215 pd=144 as=0 ps=0
M1615 a_n33822_n13887# a0 vdd w_n33912_n13914# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1616 vdd comp_b2 a_n30123_n10062# w_n29898_n10233# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1617 a_n33822_n10143# b3 a_n33822_n10269# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1618 comp_b3 a_n30330_n4554# a_n30123_n4122# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1619 a_n28773_n2844# x1 vdd w_n28890_n2754# pfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1620 a_n27072_n774# AlessB_2 vdd w_n27144_n792# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1621 carry3 a_n29637_8820# vdd w_n29718_8919# pfet w=45 l=18
+  ad=1620 pd=162 as=0 ps=0
M1622 a_n28710_45# comp_b3 vdd w_n28800_18# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1623 a_n33840_n3942# D gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1624 and_a0 a_n33822_n13887# vdd w_n33444_n13878# pfet w=54 l=18
+  ad=2916 pd=216 as=0 ps=0
M1625 AmoreB_0 a_n28773_n7173# vdd w_n28890_n7083# pfet w=54 l=18
+  ad=2430 pd=198 as=0 ps=0
M1626 a_n35820_n11565# s1_not a_n35820_n11691# Gnd nfet w=27 l=18
+  ad=972 pd=126 as=0 ps=0
M1627 and_a1 a_n33822_n13356# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1628 a_n27072_n5220# AmoreB_1 gnd Gnd nfet w=27 l=18
+  ad=0 pd=0 as=0 ps=0
M1629 comp_b2 comp_a2 a_n30123_n5067# w_n29898_n5436# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1630 a_n29853_5013# a_n30312_5085# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1631 and_oper_out0 a_n31851_n15237# gnd Gnd nfet w=27 l=18
+  ad=1458 pd=162 as=0 ps=0
M1632 a_n30312_9297# a_n30483_10044# vdd w_n30402_9270# pfet w=45 l=18
+  ad=0 pd=0 as=0 ps=0
M1633 gnd a_n29673_7947# a_n28791_7749# Gnd nfet w=54 l=18
+  ad=0 pd=0 as=0 ps=0
M1634 a_n28791_7749# a_n28998_7515# sum2 w_n28566_7578# pfet w=63 l=18
+  ad=0 pd=0 as=0 ps=0
M1635 AlessB_1 a_n28620_n1548# gnd Gnd nfet w=27 l=18
+  ad=1215 pd=144 as=0 ps=0
C0 w_n35910_n12060# vdd 0.28fF
C1 w_n35910_n12501# s0_not 0.93fF
C2 vdd a_n30312_3150# 0.60fF
C3 a_n30285_n7686# a_n28377_n7326# 0.06fF
C4 w_n33444_n12933# a_n33822_n12942# 2.17fF
C5 D1 a_n30483_5832# 0.99fF
C6 w_n28890_n2754# comp_b0 0.63fF
C7 a1 a0 0.82fF
C8 w_n28872_n792# vdd 0.28fF
C9 w_n28260_n9846# k 0.19fF
C10 AmoreB_0 a_n27072_n5220# 1.06fF
C11 vdd carry0 2.13fF
C12 a_n29673_10044# w_n28566_9675# 2.98fF
C13 a_n29673_9846# w_n29448_9675# 0.72fF
C14 comp_a1 a_n30123_n6282# 1.98fF
C15 w_n29205_n5004# comp_b2 0.66fF
C16 a_n33840_n2871# b2 0.60fF
C17 D1 a_n30690_7515# 1.06fF
C18 w_n33462_n1800# a_n33840_n1809# 2.17fF
C19 w_n29547_n4833# a_n30123_n5067# 0.66fF
C20 a1 a_n33822_n9135# 0.60fF
C21 w_n29898_n5436# a_n30123_n5265# 0.72fF
C22 w_n29898_n11250# vdd 0.48fF
C23 b3 D3 0.11fF
C24 a_n30285_n7686# a_n28773_n7173# 0.80fF
C25 w_n28737_n1458# a_n28620_n1548# 1.57fF
C26 w_n30402_5058# a_n30312_5085# 0.42fF
C27 w_n29718_2772# carry0 0.14fF
C28 gnd a_n28998_7515# 0.60fF
C29 w_n33930_n3312# b1 0.93fF
C30 w_n29934_5094# a_n29853_5013# 0.19fF
C31 b1 D2 0.12fF
C32 vdd b2 0.27fF
C33 w_n33930_n891# vdd 0.28fF
C34 comp_b2 comp_a0 0.39fF
C35 comp_b1 x1 0.86fF
C36 w_n29547_n9630# vdd 2.02fF
C37 vdd a_n30483_3897# 0.60fF
C38 adsub_b2 adsub_a1 0.67fF
C39 comp_b3 x3 0.62fF
C40 w_n29898_n2124# a_n30123_n1755# 1.20fF
C41 gnd a_n29457_n9828# 1.60fF
C42 D1 b0 0.19fF
C43 a_n30690_9612# adsub_b3 1.00fF
C44 w_n29898_n162# vdd 0.48fF
C45 a0 a_n33822_n13887# 0.60fF
C46 w_n30258_7578# adsub_b2 1.86fF
C47 w_n29898_n3420# comp_a0 2.98fF
C48 gnd a_n30330_n3483# 0.60fF
C49 w_n29547_n11943# a_n29457_n12141# 0.19fF
C50 a2 a_n33822_n8721# 0.60fF
C51 w_n28332_n4275# a_n28710_n4284# 2.17fF
C52 w_n29178_n4194# b3_not 0.19fF
C53 vdd and_a2 0.62fF
C54 w_n33912_n9162# vdd 0.28fF
C55 a_n28998_7515# sum2 0.99fF
C56 w_n33444_n12438# a_n33822_n12447# 2.17fF
C57 comp_a3 comp_a0 0.49fF
C58 w_n28566_5463# a_n29673_5832# 2.98fF
C59 w_n29448_5463# a_n29673_5634# 0.72fF
C60 w_n33912_n15849# a_n33822_n15822# 0.42fF
C61 w_n30258_3528# vdd 0.48fF
C62 w_n29898_n6453# comp_b1 2.98fF
C63 w_n33912_n9693# a0 0.93fF
C64 vdd a_n30312_7200# 0.60fF
C65 adsub_b3 adsub_a1 0.67fF
C66 w_n29898_n9288# comp_b3 2.98fF
C67 a_n29673_3897# a_n28791_3699# 1.98fF
C68 comp_a2 comp_b0 1.02fF
C69 a3 D2 0.10fF
C70 w_n31473_n14364# a_n31851_n14373# 2.17fF
C71 w_n33912_n14409# a_n33822_n14382# 0.42fF
C72 w_n29898_n7749# vdd 0.48fF
C73 sum3 w_n28566_9675# 1.20fF
C74 gnd AlessB_0 1.07fF
C75 b3 b0 0.95fF
C76 b2 b1 0.95fF
C77 vdd a_n30285_n7686# 0.02fF
C78 a_n29673_10044# sum3 1.55fF
C79 gnd a1 3.27fF
C80 w_n31473_n15228# and_oper_out0 0.19fF
C81 gnd and_b2 0.60fF
C82 w_n30258_5463# vdd 0.48fF
C83 vdd a_n30123_n1755# 1.04fF
C84 comp_a3 a_n28710_n4284# 0.60fF
C85 w_n33912_n15849# vdd 0.28fF
C86 w_n29898_n11250# comp_a1 1.86fF
C87 adsub_a1 a_n29673_5634# 3.02fF
C88 w_n29448_7578# adsub_a2 1.86fF
C89 a_n30483_7947# a_n29673_7749# 1.98fF
C90 w_n33912_n8748# a_n33822_n8721# 0.42fF
C91 w_n27576_n5085# vdd 7.49fF
C92 vdd w_n29376_9333# 0.28fF
C93 adsub_a3 a_n30312_9297# 1.81fF
C94 vdd a_n29673_3897# 1.21fF
C95 x3 comp_a0 0.41fF
C96 w_n27576_n5085# AmoreB 0.14fF
C97 vdd a_n30123_n6084# 1.04fF
C98 w_n33444_n14868# vdd 1.86fF
C99 a_n30330_n3483# a_n30123_n3051# 0.99fF
C100 w_n27144_n792# AlessB_0 1.41fF
C101 w_n29547_n3888# vdd 2.02fF
C102 vdd s1_not 0.27fF
C103 comp_b2 a_n30123_n738# 0.99fF
C104 a2 D2 0.12fF
C105 w_n33930_n1305# a_n33840_n1278# 0.42fF
C106 comp_a2 comp_b2 1.13fF
C107 w_n31941_n14796# a_n31851_n14769# 0.42fF
C108 comp_a2 a_n30330_n5499# 0.80fF
C109 w_n29898_n7749# a_n30330_n7812# 1.29fF
C110 w_n28890_n7083# a_n30285_n7686# 0.63fF
C111 a_n29565_8811# w_n29718_8919# 3.02fF
C112 a_n30330_n7812# a_n30285_n7686# 1.00fF
C113 w_n33930_n2898# b2 0.93fF
C114 w_n28566_5463# sum1 1.20fF
C115 w_n29178_n4194# comp_b3 0.66fF
C116 a3 b2 0.82fF
C117 w_n33912_n13914# vdd 0.28fF
C118 w_n35910_n12915# s0 0.93fF
C119 w_n28890_n2754# x3 0.84fF
C120 adsub_b1 a_n30483_5832# 1.16fF
C121 a_n30330_n12609# a_n30123_n12177# 0.99fF
C122 w_n33462_n3276# vdd 1.86fF
C123 vdd a_n33822_n8226# 0.60fF
C124 a_n30483_10044# a_n29673_10044# 0.99fF
C125 a_n29673_5832# a_n28791_5634# 1.98fF
C126 w_n33912_n10170# D2 0.93fF
C127 vdd a_n29565_4599# 0.60fF
C128 x2 a_n28773_n7173# 1.72fF
C129 a_n30312_9297# w_n29934_9306# 2.17fF
C130 carry2 a_n28791_9846# 1.98fF
C131 w_n29547_n11943# vdd 2.07fF
C132 comp_b0 a_n30330_n3483# 1.00fF
C133 comp_a3 comp_a2 1.99fF
C134 gnd x1 0.62fF
C135 comp_a1 a_n30285_n7686# 0.04fF
C136 w_n29898_n2124# vdd 0.48fF
C137 comp_a1 a_n30123_n1755# 1.27fF
C138 w_n28566_7578# a_n28998_7515# 1.29fF
C139 a_n30330_n225# comp_b3 0.60fF
C140 w_n29718_2772# a_n29637_2673# 0.96fF
C141 w_n33912_n8748# D2 0.93fF
C142 carry2 w_n29376_9333# 0.93fF
C143 w_n35442_n12465# a_n35820_n12474# 2.17fF
C144 gnd a_n29286_9360# 0.60fF
C145 w_n28872_n5121# b2_not 0.93fF
C146 w_n29448_5463# a_n30483_5832# 2.98fF
C147 w_n30258_5463# a_n30483_5634# 0.72fF
C148 w_n33444_n15813# and_b0 0.19fF
C149 w_n28332_54# AlessB_3 0.19fF
C150 w_n36243_n12096# vdd 0.89fF
C151 w_n33912_n14904# D3 0.93fF
C152 w_n29718_4707# a_n29565_4599# 3.02fF
C153 vdd a_n33822_n15822# 0.60fF
C154 a2 b2 0.82fF
C155 w_n27576_n756# vdd 1.86fF
C156 w_n28260_n9846# a_n28152_n9828# 1.57fF
C157 w_n33930_n891# a2 0.93fF
C158 w_n28908_3222# a_n29286_3213# 2.17fF
C159 a_n29673_10044# w_n29448_9675# 1.20fF
C160 comp_a1 a_n30123_n6084# 0.99fF
C161 w_n29898_n5436# a_n30123_n5067# 1.20fF
C162 D a1 0.07fF
C163 comp_b1 a_n30123_n11079# 0.99fF
C164 gnd D0 0.60fF
C165 a_n30330_n6516# a_n30123_n6084# 0.99fF
C166 a_n31851_n15237# and_b0 0.60fF
C167 w_n33912_n11079# vdd 0.28fF
C168 w_n35910_n11592# s0_not 0.93fF
C169 w_n28890_n7083# a_n28773_n7173# 1.57fF
C170 w_n33930_n3312# a_n33840_n3285# 0.42fF
C171 w_n29934_5094# a_n30312_5085# 2.17fF
C172 vdd a_n33840_n2871# 0.60fF
C173 w_n33462_n855# vdd 1.86fF
C174 a_n30483_5832# adsub_a1 1.55fF
C175 w_n29898_n1107# a_n30330_n1170# 1.29fF
C176 w_n28890_n2754# a_n28773_n2844# 1.57fF
C177 x3 comp_a2 0.41fF
C178 gnd a_n30330_n12609# 0.60fF
C179 vdd x2 2.76fF
C180 gnd a_n29673_10044# 1.02fF
C181 comp_b1 a_n28620_n1548# 0.80fF
C182 w_n33912_n14409# b3 0.93fF
C183 w_n33444_n11574# comp_b0 0.19fF
C184 w_n29898_n10233# vdd 0.48fF
C185 w_n33912_n10665# a_n33822_n10638# 0.42fF
C186 w_n28737_n1458# a1_not 0.63fF
C187 w_n35442_n12879# D3 0.19fF
C188 w_n29376_5121# carry0 0.93fF
C189 w_n29718_2772# vdd 2.78fF
C190 w_n30258_7578# a_n30690_7515# 1.29fF
C191 w_n29898_n3420# a_n30330_n3483# 1.29fF
C192 vdd a_n33822_n10143# 0.60fF
C193 comp_a3 a_n30123_9# 1.98fF
C194 w_n29898_n162# comp_b3 1.86fF
C195 gnd adsub_b0 1.41fF
C196 s0 a_n35820_n12888# 0.60fF
C197 adsub_a2 a_n30312_7200# 1.81fF
C198 w_n33444_n9126# vdd 1.86fF
C199 w_n29898_n2124# comp_a1 2.98fF
C200 a_n30690_3465# adsub_b0 1.00fF
C201 w_n29448_5463# a_n29673_5832# 1.20fF
C202 w_n33444_n15813# a_n33822_n15822# 2.17fF
C203 w_n29718_4707# vdd 2.78fF
C204 carry1 carry0 0.60fF
C205 w_n35442_n11556# D0 0.19fF
C206 a3 a_n33822_n8226# 0.60fF
C207 a1 b3 0.82fF
C208 w_n26901_n9846# equals_d 0.93fF
C209 temp a_n28152_n9828# 0.80fF
C210 w_n33912_n11079# b1 0.93fF
C211 gnd a_n29853_5013# 0.60fF
C212 w_n28890_n7083# x2 0.77fF
C213 w_n28890_n7083# vdd 11.51fF
C214 w_n30402_5058# adsub_b1 0.05fF
C215 D1 a_n30483_7749# 1.98fF
C216 gnd a_n29286_3213# 0.60fF
C217 w_n29718_6822# vdd 2.78fF
C218 b2 D3 0.10fF
C219 comp_b0 x1 0.41fF
C220 comp_a3 a_n30123_n4320# 1.98fF
C221 b0 D2 0.12fF
C222 a_n29565_8811# a_n29637_8820# 1.62fF
C223 vdd b1 0.27fF
C224 w_n33444_n15813# vdd 1.86fF
C225 comp_b3 a_n30285_n7686# 0.27fF
C226 w_n29448_7578# a_n29880_7515# 1.29fF
C227 adsub_a1 a_n29673_5832# 2.03fF
C228 comp_b0 a_n30123_n12375# 0.99fF
C229 a_n30483_7947# a_n29673_7947# 0.99fF
C230 vdd w_n30402_9270# 0.28fF
C231 w_n33444_n8712# a_n33822_n8721# 2.17fF
C232 w_n28404_n5085# vdd 1.75fF
C233 w_n28872_n5121# comp_a2 0.93fF
C234 a_n30330_n4554# a_n30123_n4122# 0.99fF
C235 vdd carry2 1.76fF
C236 w_n29718_6822# a_n29637_6723# 0.96fF
C237 w_n33912_n11610# D2 0.93fF
C238 x2 comp_a1 0.04fF
C239 w_n33444_n10629# comp_b2 0.19fF
C240 vdd a_n29457_n10845# 0.80fF
C241 vdd comp_a1 1.52fF
C242 gnd comp_b1 5.21fF
C243 w_n31473_n14760# vdd 1.14fF
C244 vdd a_n31851_n15237# 0.41fF
C245 D1 a_n30483_9846# 1.98fF
C246 w_n28260_n9846# a_n29457_n9828# 0.63fF
C247 w_n29376_3186# a_n29673_3897# 0.93fF
C248 w_n29898_n4491# vdd 0.48fF
C249 carry0 a_n29286_5148# 1.81fF
C250 w_n28908_7272# a_n29286_7263# 2.17fF
C251 w_n33912_n10665# D2 0.93fF
C252 gnd adsub_a0 2.13fF
C253 vdd and_a1 1.04fF
C254 vdd adsub_b2 1.22fF
C255 gnd a_n30483_7947# 0.74fF
C256 w_n33930_n2898# a_n33840_n2871# 0.42fF
C257 w_n33444_n13878# vdd 1.86fF
C258 w_n27144_n792# AlessB_3 2.24fF
C259 a_n30690_5400# a_n30483_5832# 0.99fF
C260 w_n33444_n9126# comp_a1 0.19fF
C261 comp_b0 a_n30330_n12609# 1.06fF
C262 w_n31941_n14400# and_a2 0.93fF
C263 comp_b2 x1 0.41fF
C264 w_n27144_n792# AlessB_2 0.80fF
C265 w_n28737_n5787# a_n28620_n5877# 1.57fF
C266 a_n30483_9846# w_n30258_9675# 0.72fF
C267 w_n33930_n2898# vdd 0.28fF
C268 a_n30483_10044# w_n29448_9675# 2.98fF
C269 gnd s0_not 0.46fF
C270 gnd a_n30330_n1170# 0.60fF
C271 D1 D0 0.99fF
C272 w_n33462_n1269# a_n33840_n1278# 2.17fF
C273 vdd a3 0.54fF
C274 b2 b0 0.95fF
C275 w_n30402_5058# adsub_a1 0.93fF
C276 gnd a0 3.27fF
C277 w_n29898_n12546# vdd 0.48fF
C278 w_n28737_n1458# x3 0.81fF
C279 w_n35910_n12060# s0 1.12fF
C280 w_n29718_6822# carry2 0.14fF
C281 w_n33912_n15849# D3 0.93fF
C282 gnd a_n29286_7263# 0.60fF
C283 a_n30483_10044# gnd 0.74fF
C284 adsub_b3 vdd 1.22fF
C285 w_n33930_n1836# vdd 0.28fF
C286 a_n29673_5832# carry0 0.09fF
C287 a_n30330_n2187# a_n30123_n1755# 0.99fF
C288 comp_a3 x1 0.04fF
C289 w_n30258_5463# a_n30483_5832# 1.20fF
C290 w_n28872_n5121# a_n28782_n5094# 0.42fF
C291 w_n31941_n15264# and_b0 0.93fF
C292 w_n35442_n12024# vdd 1.86fF
C293 AlessB_0 a_n27072_n891# 1.06fF
C294 w_n28404_n756# vdd 1.75fF
C295 w_n33930_n2403# D 0.93fF
C296 w_n33912_n10665# b2 0.93fF
C297 D1 adsub_b0 0.45fF
C298 w_n33444_n14373# and_b3 0.19fF
C299 w_n29934_3159# a_n29853_3078# 0.19fF
C300 w_n30402_3123# a_n30312_3150# 0.42fF
C301 w_n29898_n5436# comp_b2 3.54fF
C302 comp_b2 a_n28782_n765# 0.60fF
C303 comp_a1 a_n30330_n6516# 1.77fF
C304 w_n33462_n855# adsub_a2 0.19fF
C305 vdd a2 1.14fF
C306 comp_b1 a_n30123_n10881# 1.27fF
C307 w_n29898_n5436# a_n30330_n5499# 1.29fF
C308 gnd and_b3 0.60fF
C309 w_n33444_n11043# vdd 1.86fF
C310 comp_b2 a_n30123_n5265# 1.98fF
C311 w_n35910_n11592# a_n35820_n11565# 0.42fF
C312 w_n33912_n13914# D3 0.93fF
C313 gnd a_n29673_7947# 1.02fF
C314 vdd adsub_a2 1.81fF
C315 w_n33462_n3276# a_n33840_n3285# 2.17fF
C316 comp_b2 a_n30123_n10062# 0.99fF
C317 a_n29880_3465# adsub_a0 1.05fF
C318 a3 b1 0.82fF
C319 w_n33930_n1305# D 0.93fF
C320 w_n33930_n396# vdd 0.28fF
C321 a_n30483_5832# a_n29880_5400# 1.60fF
C322 D1 a_n29286_3213# 1.81fF
C323 comp_b0 comp_b1 0.98fF
C324 w_n33444_n10629# a_n33822_n10638# 2.17fF
C325 w_n33912_n10170# vdd 0.28fF
C326 x3 x1 0.27fF
C327 w_n33912_n15849# b0 0.93fF
C328 comp_b3 x2 0.41fF
C329 w_n27576_n5085# AmoreB_0 1.41fF
C330 vdd comp_b3 2.00fF
C331 vdd and_b1 1.06fF
C332 w_n29376_3186# vdd 0.28fF
C333 comp_b0 a_n30123_n3249# 1.98fF
C334 w_n30402_3123# a_n30483_3897# 0.93fF
C335 adsub_b3 w_n30402_9270# 0.05fF
C336 adsub_a3 vdd 1.81fF
C337 carry0 sum1 0.99fF
C338 a_n29673_7947# sum2 1.55fF
C339 comp_a3 a_n30123_207# 1.27fF
C340 gnd a_n30690_3465# 0.60fF
C341 w_n29898_n2124# a_n30330_n2187# 1.29fF
C342 w_n33912_n8748# vdd 0.28fF
C343 w_n33912_n10170# a_n33822_n10143# 0.42fF
C344 vdd a_n29565_8811# 0.60fF
C345 w_n33930_n2403# b3 0.93fF
C346 w_n28044_n5121# a_n27954_n5094# 0.42fF
C347 w_n29376_5121# vdd 0.28fF
C348 AmoreB_3 a_n27072_n5220# 1.04fF
C349 w_n28872_n792# a2_not 0.93fF
C350 comp_a3 a_n30123_n9117# 1.98fF
C351 a2 b1 0.82fF
C352 a_n33840_n1809# a0 0.60fF
C353 w_n34488_n1134# D0 0.80fF
C354 a_n29457_n12141# a_n28152_n9828# 0.80fF
C355 gnd a_n30330_n4554# 0.60fF
C356 D1 adsub_a0 0.07fF
C357 w_n33444_n14373# a_n33822_n14382# 2.17fF
C358 w_n29214_n5850# vdd 1.29fF
C359 a1 D2 0.12fF
C360 D1 a_n30483_7947# 0.99fF
C361 vdd a_n33822_n11583# 0.60fF
C362 comp_a2 a_n30285_n7686# 0.27fF
C363 D a0 0.07fF
C364 w_n29376_7236# vdd 0.28fF
C365 comp_a3 a_n30123_n4122# 0.99fF
C366 vdd carry1 1.27fF
C367 comp_b2 comp_b1 2.24fF
C368 vdd a_n33840_n3285# 0.60fF
C369 w_n31941_n15264# vdd 0.28fF
C370 w_n29898_n1107# comp_b2 1.86fF
C371 vdd a_n28710_45# 0.41fF
C372 a_n29880_5400# a_n29673_5832# 0.99fF
C373 comp_b0 a_n30123_n12177# 1.27fF
C374 gnd and_a3 0.66fF
C375 a_n29565_2664# a_n29637_2673# 1.62fF
C376 vdd w_n29934_9306# 1.86fF
C377 w_n29205_n5004# vdd 1.92fF
C378 s1_not s0 0.04fF
C379 w_n29268_n7146# b0_not 0.19fF
C380 x3 a_n28224_n1701# 0.06fF
C381 vdd a_n26811_n9819# 0.41fF
C382 x1 a_n28773_n2844# 1.58fF
C383 vdd a_n33822_n15291# 0.60fF
C384 w_n31941_n14400# vdd 0.28fF
C385 D1 a_n30483_10044# 0.99fF
C386 x2 comp_a0 0.41fF
C387 w_n30258_7578# a_n30483_7749# 0.72fF
C388 w_n29547_n9630# a_n29457_n9828# 0.19fF
C389 w_n29547_n2817# a_n30123_n3051# 0.66fF
C390 w_n29898_n3420# a_n30123_n3249# 0.72fF
C391 vdd comp_a0 0.96fF
C392 vdd a_n30483_5832# 0.60fF
C393 adsub_a3 w_n30402_9270# 0.93fF
C394 w_n28566_3528# sum0 1.20fF
C395 w_n33930_n3843# vdd 0.28fF
C396 comp_a3 comp_b1 0.65fF
C397 comp_b3 comp_a1 1.61fF
C398 w_n29718_4707# carry1 0.14fF
C399 w_n30402_7173# a_n30312_7200# 0.42fF
C400 w_n29934_7209# a_n29853_7128# 0.19fF
C401 a3 a2 0.82fF
C402 a_n30330_n1170# comp_b2 0.60fF
C403 w_n28332_n4275# AmoreB_3 0.19fF
C404 gnd a_n29880_3465# 0.60fF
C405 vdd a_n33822_n13356# 0.60fF
C406 w_n29898_n162# a_n30123_9# 0.72fF
C407 w_n29547_441# a_n30123_207# 0.66fF
C408 w_n33912_n14904# a_n33822_n14877# 0.42fF
C409 carry1 a_n28791_7749# 1.98fF
C410 w_n33444_n12438# and_a3 0.19fF
C411 adsub_b0 a_n30483_3699# 1.98fF
C412 b0 a_n33822_n15822# 0.60fF
C413 w_n29898_n4491# comp_b3 2.98fF
C414 w_n33912_n13383# vdd 0.28fF
C415 w_n33930_n396# a3 0.93fF
C416 and_a1 and_b1 2.13fF
C417 a_n30483_10044# w_n30258_9675# 1.20fF
C418 w_n28890_n2754# x2 0.77fF
C419 a0 b3 0.82fF
C420 w_n28890_n2754# vdd 11.51fF
C421 a1 b2 0.82fF
C422 vdd a_n28710_n4284# 0.41fF
C423 w_n31473_n14364# and_oper_out2 0.19fF
C424 D1 sum0 0.99fF
C425 vdd a_n29286_5148# 0.60fF
C426 w_n33912_n9693# D2 0.93fF
C427 adsub_b3 adsub_a2 0.41fF
C428 a_n33840_n3285# b1 0.60fF
C429 w_n36243_n12096# s0 0.66fF
C430 w_n33912_n12474# vdd 0.28fF
C431 vdd a_n29565_2664# 0.60fF
C432 w_n29547_n8685# a_n30123_n8919# 0.66fF
C433 b1 D3 0.13fF
C434 w_n29898_n9288# a_n30123_n9117# 0.72fF
C435 a_n31851_n13896# and_b3 0.60fF
C436 a_n28998_3465# sum0 0.99fF
C437 carry2 carry1 0.60fF
C438 vdd b0 0.27fF
C439 gnd comp_b0 4.26fF
C440 w_n28737_n5787# b1_not 0.63fF
C441 w_n29898_n6453# a_n30123_n6282# 0.72fF
C442 w_n29547_n5850# a_n30123_n6084# 0.66fF
C443 w_n33462_n1800# vdd 1.86fF
C444 a_n29673_5832# a_n28998_5400# 1.08fF
C445 gnd D 5.33fF
C446 w_n29448_7578# a_n29673_7749# 0.72fF
C447 w_n28566_7578# a_n29673_7947# 2.98fF
C448 w_n33912_n8253# D2 0.93fF
C449 x3 a_n27954_n5094# 1.21fF
C450 w_n29718_2772# a_n29565_2664# 3.02fF
C451 x3 comp_b1 0.04fF
C452 a_n28998_9612# carry2 2.85fF
C453 gnd a_n29853_9225# 0.60fF
C454 b1 a_n33822_n15291# 0.60fF
C455 w_n31941_n15264# a_n31851_n15237# 0.42fF
C456 w_n33912_n11610# vdd 0.28fF
C457 w_n29547_n1521# x1 0.19fF
C458 w_n33912_n9162# a1 0.93fF
C459 and_a2 and_b2 0.87fF
C460 w_n33444_n8217# comp_a3 0.19fF
C461 w_n29205_n675# vdd 1.92fF
C462 D1 gnd 8.91fF
C463 w_n29547_n2817# x0 0.19fF
C464 a_n30330_n2187# comp_a1 1.73fF
C465 w_n31941_n13923# and_b3 0.93fF
C466 D1 a_n30690_3465# 1.03fF
C467 vdd a_n29673_5832# 1.21fF
C468 w_n29934_3159# a_n30312_3150# 2.17fF
C469 AlessB_3 a_n27072_n891# 1.04fF
C470 vdd s0 0.60fF
C471 comp_a1 comp_a0 0.35fF
C472 comp_b1 a_n30330_n11313# 0.99fF
C473 gnd a_n28998_3465# 0.60fF
C474 vdd and_a0 0.77fF
C475 comp_b2 a_n30123_n5067# 1.27fF
C476 w_n35442_n11556# a_n35820_n11565# 2.17fF
C477 w_n33912_n10665# vdd 0.28fF
C478 a_n30330_n5499# a_n30123_n5067# 0.99fF
C479 comp_b2 a_n30123_n9864# 1.27fF
C480 w_n28890_n7083# AmoreB_0 0.19fF
C481 w_n33462_n360# vdd 1.86fF
C482 a_n30330_n10296# a_n30123_n9864# 0.99fF
C483 a3 D3 0.04fF
C484 vdd a_n35820_n12474# 0.60fF
C485 vdd a_n30123_n738# 1.04fF
C486 w_n28737_n1458# AlessB_1 0.19fF
C487 comp_a2 x2 0.92fF
C488 adsub_b1 adsub_a0 0.41fF
C489 b2 a_n33822_n14877# 0.60fF
C490 gnd comp_b2 5.33fF
C491 vdd comp_a2 1.86fF
C492 gnd a_n30330_n5499# 0.60fF
C493 w_n33444_n10134# vdd 1.86fF
C494 gnd a_n30330_n10296# 0.60fF
C495 w_n33912_n8748# a2 0.93fF
C496 w_n29898_n10233# comp_a2 1.86fF
C497 x3 a_n28620_n1548# 1.67fF
C498 b1 b0 0.95fF
C499 gnd b3 3.49fF
C500 w_n28800_n4311# comp_a3 0.93fF
C501 w_n30402_3123# vdd 0.28fF
C502 vdd a_n31851_n14769# 0.41fF
C503 comp_b0 a_n30123_n3051# 0.99fF
C504 w_n29448_3528# adsub_a0 1.86fF
C505 a_n30690_7515# adsub_b2 1.00fF
C506 vdd a_n29565_6714# 0.60fF
C507 vdd a_n33822_n9666# 0.60fF
C508 a_n28998_5400# sum1 0.99fF
C509 comp_b1 a_n30123_n1953# 1.98fF
C510 w_n28566_7578# sum2 1.20fF
C511 w_n33444_n14868# and_b2 0.19fF
C512 vdd a_n33822_n12942# 0.60fF
C513 a_n30330_n225# a_n30123_207# 0.99fF
C514 w_n33444_n8712# vdd 1.86fF
C515 w_n33444_n10134# a_n33822_n10143# 2.17fF
C516 gnd a_n30330_n9351# 0.60fF
C517 w_n29898_n12546# comp_a0 1.86fF
C518 w_n33930_n2403# a_n33840_n2376# 0.42fF
C519 w_n27576_n5085# AmoreB_2 0.99fF
C520 w_n28044_n5121# a_n28323_n5166# 0.93fF
C521 x3 a_n28620_n5877# 1.67fF
C522 a_n29565_6714# a_n29637_6723# 1.62fF
C523 w_n30402_5058# vdd 0.28fF
C524 gnd comp_a3 5.43fF
C525 a_n30330_n9351# a_n30123_n8919# 0.99fF
C526 w_n28872_n792# a_n28782_n765# 0.42fF
C527 x2 a_n28494_n6030# 0.06fF
C528 w_n28737_n5787# x3 0.81fF
C529 comp_a3 a_n30123_n8919# 0.99fF
C530 b3 a_n33822_n14382# 0.60fF
C531 a_n29457_n10845# a_n28152_n9828# 0.80fF
C532 a2 D3 0.10fF
C533 w_n29547_n5850# vdd 1.95fF
C534 comp_b1 a_n30123_n6282# 1.98fF
C535 w_n30402_7173# vdd 0.28fF
C536 gnd a_n29853_3078# 0.60fF
C537 w_n33912_n12474# a3 0.93fF
C538 w_n31941_n13923# and_a3 0.93fF
C539 adsub_a0 a_n29673_3699# 3.02fF
C540 w_n33912_n15318# vdd 0.28fF
C541 a3 b0 0.82fF
C542 a_n30483_5832# a_n29673_5634# 1.98fF
C543 w_n29448_7578# a_n30483_7947# 2.98fF
C544 vdd a_n33822_n12447# 0.60fF
C545 w_n29268_n7146# comp_b0 0.66fF
C546 w_n29547_n4833# x2 0.19fF
C547 w_n29547_n4833# vdd 2.02fF
C548 vdd w_n28908_9369# 1.86fF
C549 comp_b0 a_n30123_n7578# 1.98fF
C550 s1_not a_n35820_n11691# 0.06fF
C551 w_n29718_6822# a_n29565_6714# 3.02fF
C552 comp_b1 a_n28620_n1701# 0.10fF
C553 vdd a_n28782_n5094# 1.02fF
C554 w_n28566_3528# D1 1.95fF
C555 comp_b3 a_n28710_45# 0.60fF
C556 vdd a_n29457_n9828# 0.80fF
C557 comp_a2 comp_a1 1.33fF
C558 a_n30690_9612# a_n30483_10044# 0.99fF
C559 w_n33912_n14409# vdd 0.28fF
C560 gnd x3 1.85fF
C561 w_n30258_7578# a_n30483_7947# 1.20fF
C562 s1_not a_n35820_n12159# 0.06fF
C563 w_n29898_n3420# a_n30123_n3051# 1.20fF
C564 w_n33444_n13878# and_a0 0.19fF
C565 w_n28566_3528# a_n28998_3465# 1.29fF
C566 w_n33912_n13914# a_n33822_n13887# 0.42fF
C567 w_n33462_n3807# vdd 1.86fF
C568 w_n29934_7209# a_n30312_7200# 2.17fF
C569 w_n29898_n162# a_n30123_207# 1.20fF
C570 w_n33444_n14868# a_n33822_n14877# 2.17fF
C571 w_n31473_n14760# a_n31851_n14769# 2.17fF
C572 a_n29286_9360# w_n29376_9333# 0.42fF
C573 adsub_b0 a_n30483_3897# 0.99fF
C574 w_n33462_n2862# a_n33840_n2871# 2.17fF
C575 comp_b3 comp_a0 0.68fF
C576 w_n28737_n5787# AmoreB_1 0.19fF
C577 w_n33444_n13347# vdd 1.86fF
C578 gnd a_n30330_n11313# 0.60fF
C579 gnd adsub_b1 1.72fF
C580 w_n28044_n792# a_n27954_n765# 0.42fF
C581 comp_b2 comp_b0 1.66fF
C582 a2 b0 0.82fF
C583 w_n33462_n2862# vdd 1.86fF
C584 w_n29376_7236# carry1 0.93fF
C585 D1 a_n28998_3465# 2.85fF
C586 w_n29178_135# comp_a3 0.66fF
C587 a_n28791_9846# w_n28566_9675# 0.72fF
C588 a_n29673_10044# a_n28791_9846# 1.98fF
C589 a0 D2 0.12fF
C590 vdd a1 0.27fF
C591 w_n33912_n15318# b1 0.93fF
C592 vdd and_b2 1.80fF
C593 D b3 0.09fF
C594 w_n35910_n12501# vdd 0.28fF
C595 w_n29898_n9288# a_n30123_n8919# 1.20fF
C596 adsub_a0 a_n30312_3150# 1.81fF
C597 w_n30258_3528# adsub_b0 1.86fF
C598 gnd a_n29853_7128# 0.60fF
C599 w_n29898_n3420# comp_b0 1.86fF
C600 w_n29898_n6453# a_n30123_n6084# 1.20fF
C601 w_n28737_n1458# x2 0.84fF
C602 D1 w_n30258_9675# 2.98fF
C603 vdd a_n33840_n3816# 0.60fF
C604 w_n28737_n1458# vdd 11.51fF
C605 w_n29898_n11250# comp_b1 2.98fF
C606 x3 a_n27954_n765# 1.21fF
C607 w_n29448_7578# a_n29673_7947# 1.20fF
C608 w_n33912_n8253# a_n33822_n8226# 0.42fF
C609 x1 a_n28773_n7173# 1.58fF
C610 x3 a_n28323_n5166# 0.06fF
C611 a_n29673_10044# w_n29376_9333# 0.93fF
C612 comp_a3 comp_b0 0.48fF
C613 w_n28404_n5085# a_n28782_n5094# 2.17fF
C614 w_n29205_n5004# b2_not 0.19fF
C615 gnd AmoreB_1 1.07fF
C616 w_n33444_n11574# vdd 1.86fF
C617 w_n29376_5121# a_n29286_5148# 0.42fF
C618 w_n29547_n504# x2 0.19fF
C619 a_n30690_9612# gnd 0.60fF
C620 w_n29547_n504# vdd 2.02fF
C621 w_n30402_7173# adsub_b2 0.05fF
C622 comp_b0 a_n28377_n2997# 0.06fF
C623 w_n31941_n13923# a_n31851_n13896# 0.42fF
C624 a_n29880_7515# adsub_a2 1.03fF
C625 w_n27144_n792# a_n27072_n891# 0.96fF
C626 w_n29547_n10647# a_n30123_n10881# 0.66fF
C627 w_n29898_n11250# a_n30123_n11079# 0.72fF
C628 vdd a_n33822_n13887# 0.60fF
C629 comp_b2 a_n30330_n5499# 1.73fF
C630 w_n33444_n10629# vdd 1.86fF
C631 w_n29214_n1521# a1_not 0.19fF
C632 comp_b2 a_n30330_n10296# 1.06fF
C633 w_n33912_n13383# D3 0.93fF
C634 a_n30483_3897# adsub_a0 1.55fF
C635 w_n28566_5463# a_n28791_5634# 0.72fF
C636 a_n35820_n12474# s1 0.60fF
C637 w_n28800_18# vdd 0.28fF
C638 and_a0 and_b1 0.54fF
C639 gnd adsub_a1 2.41fF
C640 a3 a_n33822_n12447# 0.60fF
C641 b0 a_n33822_n11583# 0.60fF
C642 comp_a2 a_n30123_n936# 1.98fF
C643 a1 b1 0.82fF
C644 a0 b2 0.82fF
C645 a2 a_n33822_n12942# 0.60fF
C646 w_n33912_n9693# vdd 0.28fF
C647 w_n33912_n12474# D3 0.93fF
C648 w_n29376_5121# a_n29673_5832# 0.93fF
C649 x3 comp_b0 0.41fF
C650 a_n30330_n11313# a_n30123_n10881# 0.99fF
C651 vdd a_n33822_n14877# 0.60fF
C652 w_n33462_n360# adsub_a3 0.19fF
C653 w_n34488_n1134# D 0.14fF
C654 w_n29934_3159# vdd 1.86fF
C655 w_n33912_n11610# a_n33822_n11583# 0.42fF
C656 comp_b3 comp_a2 1.33fF
C657 x2 x1 0.27fF
C658 b0 D3 0.06fF
C659 comp_a3 comp_b2 0.34fF
C660 w_n33912_n13383# a_n33822_n13356# 0.42fF
C661 comp_b1 a_n30285_n7686# 0.06fF
C662 w_n33444_n13347# and_a1 0.19fF
C663 vdd x1 1.23fF
C664 w_n29448_3528# a_n29880_3465# 1.29fF
C665 w_n33444_n10134# comp_b3 0.19fF
C666 gnd D2 4.84fF
C667 adsub_a1 a_n30312_5085# 1.81fF
C668 comp_b1 a_n30123_n1755# 0.99fF
C669 w_n29547_n3888# a_n30123_n4122# 0.66fF
C670 w_n29898_n4491# a_n30123_n4320# 0.72fF
C671 a_n31851_n14769# and_b1 0.60fF
C672 w_n33912_n8253# vdd 0.28fF
C673 w_n33462_n2862# adsub_b2 0.19fF
C674 w_n33462_n2367# a_n33840_n2376# 2.17fF
C675 vdd a_n29286_9360# 0.60fF
C676 w_n27576_n5085# a_n27954_n5094# 2.17fF
C677 gnd a_n30330_n225# 0.60fF
C678 w_n34488_n1134# D1 0.80fF
C679 w_n29934_5094# vdd 1.86fF
C680 w_n36234_n12420# s1_not 0.19fF
C681 w_n33912_n11079# a_n33822_n11052# 0.42fF
C682 and_a1 and_b2 0.54fF
C683 w_n33930_n3843# b0 0.93fF
C684 w_n28044_n5121# x3 2.64fF
C685 a_n29880_9612# adsub_a3 1.03fF
C686 w_n30402_7173# adsub_a2 0.93fF
C687 w_n33930_n891# a_n33840_n864# 0.42fF
C688 w_n31941_n15264# and_a0 0.93fF
C689 D1 a_n30483_3699# 1.98fF
C690 w_n33912_n9162# a_n33822_n9135# 0.42fF
C691 comp_b1 a_n30123_n6084# 1.27fF
C692 w_n29898_n6453# vdd 0.48fF
C693 vdd a_n33822_n11052# 0.60fF
C694 vdd D0 1.04fF
C695 a3 a1 0.82fF
C696 w_n35910_n11592# s1_not 0.93fF
C697 w_n28800_18# a3_not 0.93fF
C698 w_n29934_7209# vdd 1.86fF
C699 D1 adsub_b1 0.11fF
C700 w_n33462_n1269# adsub_a1 0.19fF
C701 adsub_a0 a_n29673_3897# 2.03fF
C702 w_n33444_n15282# vdd 1.86fF
C703 w_n28890_n7083# x1 0.74fF
C704 a_n30483_5832# a_n29673_5832# 0.99fF
C705 x3 comp_b2 0.04fF
C706 gnd carry0 1.21fF
C707 AmoreB_1 a_n27072_n5220# 1.06fF
C708 comp_b0 a_n30123_n7380# 1.27fF
C709 vdd w_n28566_9675# 0.48fF
C710 w_n29898_n5436# vdd 0.48fF
C711 vdd a_n28782_n765# 1.02fF
C712 vdd a_n29673_10044# 1.21fF
C713 w_n27576_n5085# AmoreB_3 2.24fF
C714 w_n28737_n1458# temp_less 0.63fF
C715 and_a2 and_b3 0.54fF
C716 gnd b2 3.55fF
C717 w_n29547_n9630# a_n30123_n9864# 0.66fF
C718 w_n31473_n14364# vdd 1.14fF
C719 w_n29898_n10233# a_n30123_n10062# 0.72fF
C720 vdd a_n30123_207# 1.04fF
C721 comp_b0 a_n28773_n2844# 0.80fF
C722 comp_a2 comp_a0 15.88fF
C723 w_n33444_n13878# a_n33822_n13887# 2.17fF
C724 adsub_b2 a_n30483_7749# 1.98fF
C725 w_n29268_n2817# vdd 1.62fF
C726 s0_not s1_not 4.35fF
C727 adsub_a3 a_n29673_9846# 2.83fF
C728 comp_a1 x1 1.23fF
C729 w_n33912_n11610# b0 0.93fF
C730 vdd adsub_b0 0.76fF
C731 gnd a_n30483_3897# 0.74fF
C732 comp_a3 x3 0.99fF
C733 comp_b3 a_n30123_9# 1.98fF
C734 a_n29565_8811# w_n28908_9369# 0.19fF
C735 w_n29898_n2124# comp_b1 1.86fF
C736 a_n29853_9225# w_n29718_8919# 0.80fF
C737 a_n30690_3465# a_n30483_3897# 0.99fF
C738 carry2 a_n29286_9360# 1.81fF
C739 a_n30690_9612# D1 1.06fF
C740 a2 a1 0.82fF
C741 w_n29547_n8685# a_n29457_n8883# 0.19fF
C742 w_n33912_n12969# vdd 0.28fF
C743 gnd a_n30690_5400# 0.60fF
C744 w_n27576_n756# AlessB_2 0.19fF
C745 b1 a_n33822_n11052# 0.60fF
C746 w_n28044_n792# a_n28323_n837# 0.93fF
C747 w_n33930_n2403# vdd 0.28fF
C748 w_n33912_n13914# a0 0.93fF
C749 gnd and_a2 0.60fF
C750 vdd a_n30123_n4122# 1.04fF
C751 a_n28998_7515# carry1 2.85fF
C752 w_n35910_n12501# s1 0.93fF
C753 comp_a1 a_n28620_n6030# 0.10fF
C754 w_n30402_5058# a_n30483_5832# 0.93fF
C755 vdd a_n33840_n1278# 0.60fF
C756 w_n28044_n792# x3 2.64fF
C757 vdd a_n31851_n14373# 0.41fF
C758 w_n29898_n9288# a_n30330_n9351# 1.29fF
C759 w_n36234_n12420# vdd 2.50fF
C760 vdd a_n29286_3213# 0.60fF
C761 w_n29898_n6453# comp_a1 1.86fF
C762 w_n33912_n15318# D3 0.93fF
C763 w_n33444_n12933# and_a2 0.19fF
C764 comp_b3 a_n30123_n4320# 1.98fF
C765 D1 adsub_a1 0.12fF
C766 a_n29673_3897# sum0 1.55fF
C767 w_n30258_3528# a_n30690_3465# 1.29fF
C768 w_n29898_n6453# a_n30330_n6516# 1.29fF
C769 w_n29898_n9288# comp_a3 1.86fF
C770 a_n30690_9612# w_n30258_9675# 1.29fF
C771 w_n33930_n1305# vdd 0.28fF
C772 w_n33930_n3312# D 0.93fF
C773 x3 a_n28323_n837# 0.06fF
C774 vdd AlessB_3 0.60fF
C775 w_n33444_n8217# a_n33822_n8226# 2.17fF
C776 w_n30258_7578# D1 2.98fF
C777 w_n33912_n8253# a3 0.93fF
C778 carry2 w_n28566_9675# 1.95fF
C779 gnd AlessB_1 1.07fF
C780 a_n29673_10044# carry2 0.09fF
C781 gnd a_n30285_n7686# 1.49fF
C782 vdd a_n27954_n5094# 0.60fF
C783 w_n36243_n12096# s0_not 0.19fF
C784 w_n33912_n15318# a_n33822_n15291# 0.42fF
C785 w_n35910_n11592# vdd 0.28fF
C786 x2 comp_b1 0.04fF
C787 vdd comp_b1 2.71fF
C788 w_n35910_n12915# a_n35820_n12888# 0.42fF
C789 w_n29547_n11943# a_n30123_n12177# 0.66fF
C790 w_n29898_n12546# a_n30123_n12375# 0.72fF
C791 w_n33912_n14409# D3 0.93fF
C792 w_n28908_5157# a_n29565_4599# 0.19fF
C793 w_n29718_4707# a_n29853_5013# 0.80fF
C794 w_n29898_n1107# vdd 0.48fF
C795 adsub_b3 a_n30483_9846# 1.98fF
C796 w_n29205_n675# comp_a2 0.66fF
C797 w_n31473_n13887# a_n31851_n13896# 2.17fF
C798 w_n29898_n11250# a_n30123_n10881# 1.20fF
C799 a3 D0 0.06fF
C800 gnd a_n29673_3897# 1.02fF
C801 vdd adsub_a0 1.81fF
C802 w_n29547_441# x3 0.19fF
C803 w_n26901_n9846# vdd 0.28fF
C804 gnd a_n29457_n12141# 0.80fF
C805 vdd a_n30483_7947# 0.60fF
C806 a_n30483_3897# a_n29880_3465# 1.60fF
C807 a_n30330_n3483# comp_a0 1.73fF
C808 gnd and_b0 1.20fF
C809 w_n28332_54# vdd 1.14fF
C810 gnd a_n29880_5400# 0.60fF
C811 w_n27144_n792# AlessB_1 0.99fF
C812 comp_a2 a_n30123_n738# 1.27fF
C813 a_n33840_n2376# b3 0.60fF
C814 vdd s0_not 0.73fF
C815 gnd s1_not 1.35fF
C816 D1 a_n34407_n1233# 0.60fF
C817 vdd AmoreB_3 0.60fF
C818 a1 D3 0.10fF
C819 w_n28800_18# comp_b3 0.93fF
C820 w_n33444_n9657# vdd 1.86fF
C821 w_n33912_n12474# a_n33822_n12447# 0.42fF
C822 w_n29898_n12546# a_n30330_n12609# 1.29fF
C823 w_n28566_5463# carry0 1.95fF
C824 b3 D2 0.12fF
C825 vdd a0 0.27fF
C826 D b2 0.12fF
C827 w_n35910_n12060# a_n35820_n12033# 0.42fF
C828 w_n33444_n11574# a_n33822_n11583# 2.17fF
C829 w_n33930_n891# D 0.93fF
C830 w_n28908_3222# vdd 1.86fF
C831 x2 a_n28620_n1548# 1.16fF
C832 D1 carry0 0.46fF
C833 w_n33444_n13347# a_n33822_n13356# 2.17fF
C834 vdd a_n29286_7263# 0.60fF
C835 vdd a_n33822_n9135# 0.60fF
C836 a_n30483_10044# vdd 0.60fF
C837 a_n29673_5832# sum1 1.55fF
C838 w_n29898_n4491# a_n30123_n4122# 1.20fF
C839 w_n31941_n14400# and_b2 0.93fF
C840 vdd a_n30123_n12177# 1.04fF
C841 w_n33444_n8217# vdd 1.86fF
C842 comp_b3 x1 0.41fF
C843 w_n33444_n8712# comp_a2 0.19fF
C844 carry2 sum3 0.99fF
C845 a2 D0 0.06fF
C846 w_n33444_n11043# a_n33822_n11052# 2.17fF
C847 w_n28908_5157# vdd 1.86fF
C848 a1 a_n33822_n13356# 0.60fF
C849 x3 a_n28773_n2844# 1.16fF
C850 w_n33930_n3843# a_n33840_n3816# 0.42fF
C851 x2 a_n28620_n5877# 1.16fF
C852 w_n28404_n756# a_n28782_n765# 2.17fF
C853 w_n29205_n675# a2_not 0.19fF
C854 w_n33462_n855# a_n33840_n864# 2.17fF
C855 w_n28872_n792# comp_b2 0.93fF
C856 a_n29457_n9828# a_n28152_n9828# 0.80fF
C857 w_n33912_n13383# a1 0.93fF
C858 comp_a1 comp_b1 0.80fF
C859 a_n30330_n225# comp_a3 1.80fF
C860 D1 a_n30483_3897# 0.99fF
C861 adsub_a2 a_n29673_7749# 2.83fF
C862 w_n33444_n9126# a_n33822_n9135# 2.17fF
C863 w_n28737_n5787# x2 0.84fF
C864 comp_b1 a_n30330_n6516# 1.73fF
C865 w_n28737_n5787# vdd 11.51fF
C866 w_n28890_n2754# AlessB_0 0.19fF
C867 vdd a_n33840_n864# 0.60fF
C868 w_n35442_n12465# D2 0.19fF
C869 vdd and_b3 1.06fF
C870 w_n28800_18# a_n28710_45# 0.42fF
C871 w_n28908_7272# vdd 1.86fF
C872 D1 a_n30690_5400# 1.06fF
C873 vdd a_n29673_7947# 1.21fF
C874 a_n29880_3465# a_n29673_3897# 0.99fF
C875 w_n31473_n15228# vdd 1.14fF
C876 w_n28260_n9846# temp 0.63fF
C877 gnd a_n28998_5400# 0.60fF
C878 w_n29898_n7749# comp_b0 2.98fF
C879 comp_b0 a_n30285_n7686# 0.75fF
C880 w_n28800_n4311# vdd 0.28fF
C881 vdd w_n29448_9675# 0.48fF
C882 a0 b1 0.82fF
C883 a1 b0 0.82fF
C884 b3 b2 1.08fF
C885 comp_a1 a_n30123_n11079# 1.98fF
C886 w_n33444_n15282# and_b1 0.19fF
C887 vdd a_n30123_n5067# 1.04fF
C888 comp_a2 a_n28782_n5094# 0.60fF
C889 w_n30258_3528# D1 2.98fF
C890 w_n29898_n7749# a_n30123_n7578# 0.72fF
C891 w_n28890_n7083# b0_not 0.63fF
C892 carry3 w_n29718_8919# 0.14fF
C893 w_n29547_n7146# a_n30123_n7380# 0.66fF
C894 a_n30285_n7686# a_n30123_n7578# 1.98fF
C895 vdd a_n30123_n9864# 1.04fF
C896 a_n33840_n3816# b0 0.60fF
C897 w_n27576_n5085# a_n27072_n5220# 0.96fF
C898 w_n33444_n14373# vdd 1.86fF
C899 w_n29898_n10233# a_n30123_n9864# 1.20fF
C900 vdd a_n33840_n369# 0.60fF
C901 adsub_b2 adsub_a0 0.41fF
C902 w_n28260_n9846# a_n29457_n8883# 0.63fF
C903 w_n33912_n12969# a2 0.93fF
C904 w_n28890_n2754# a0_not 0.63fF
C905 w_n29448_3528# a_n29673_3699# 0.72fF
C906 w_n28566_3528# a_n29673_3897# 2.98fF
C907 adsub_b2 a_n30483_7947# 1.16fF
C908 a_n30483_10044# w_n30402_9270# 0.93fF
C909 gnd x2 1.31fF
C910 gnd vdd 14.95fF
C911 adsub_a3 a_n29673_10044# 1.84fF
C912 a_n35820_n11565# s1_not 0.60fF
C913 w_n29547_n2817# vdd 1.95fF
C914 carry0 a_n28791_5634# 1.98fF
C915 w_n30258_5463# D1 2.98fF
C916 a_n29673_7947# a_n28791_7749# 1.98fF
C917 comp_b3 a_n30123_207# 0.99fF
C918 vdd a_n30123_n8919# 1.04fF
C919 x1 comp_a0 0.41fF
C920 w_n33444_n12933# vdd 1.86fF
C921 and_a0 and_b2 0.54fF
C922 w_n27576_n756# a_n27954_n765# 2.17fF
C923 comp_b3 a_n30123_n9117# 0.99fF
C924 comp_a0 a_n30123_n12375# 1.98fF
C925 w_n33462_n2367# vdd 1.86fF
C926 w_n26433_n9810# AequalsB 0.19fF
C927 w_n34488_n1134# a_n34407_n1233# 0.96fF
C928 w_n29898_n162# comp_a3 2.98fF
C929 adsub_b3 adsub_a0 0.41fF
C930 D1 a_n29673_3897# 0.09fF
C931 vdd a_n30312_5085# 0.60fF
C932 w_n35910_n12501# a_n35820_n12474# 0.42fF
C933 comp_a1 a_n28620_n5877# 0.80fF
C934 w_n36234_n12420# s1 0.66fF
C935 comp_b2 a_n30285_n7686# 0.27fF
C936 w_n29448_5463# adsub_a1 1.86fF
C937 a3 a0 0.82fF
C938 vdd a_n33822_n14382# 0.60fF
C939 w_n28737_n5787# comp_a1 0.63fF
C940 w_n33444_n12438# vdd 1.86fF
C941 w_n28890_n2754# x1 0.74fF
C942 comp_b3 a_n30123_n4122# 1.27fF
C943 a_n29673_3897# a_n28998_3465# 1.08fF
C944 w_n26901_n9846# k 0.93fF
C945 w_n27144_n792# vdd 3.84fF
C946 w_n33444_n11043# comp_b1 0.19fF
C947 w_n29376_3186# a_n29286_3213# 0.42fF
C948 vdd and_a3 0.62fF
C949 vdd a_n27954_n765# 0.60fF
C950 a_n28998_9612# w_n28566_9675# 1.29fF
C951 s1_not a_n35820_n12033# 0.60fF
C952 gnd a_n30330_n7812# 0.60fF
C953 a_n29673_10044# a_n28998_9612# 1.08fF
C954 w_n33930_n1836# a0 0.93fF
C955 temp_less a_n28620_n1548# 0.80fF
C956 w_n33444_n15282# a_n33822_n15291# 2.17fF
C957 w_n31473_n15228# a_n31851_n15237# 2.17fF
C958 w_n29547_n7146# a_n29457_n7344# 0.19fF
C959 w_n35442_n11556# vdd 1.86fF
C960 and_a1 and_b3 0.54fF
C961 w_n29898_n12546# a_n30123_n12177# 1.20fF
C962 w_n35442_n12879# a_n35820_n12888# 2.17fF
C963 w_n29898_n1107# a_n30123_n936# 0.72fF
C964 gnd b1 3.57fF
C965 w_n29547_n504# a_n30123_n738# 0.66fF
C966 adsub_b3 a_n30483_10044# 1.16fF
C967 w_n33462_n1269# vdd 1.86fF
C968 comp_a3 a_n30285_n7686# 0.01fF
C969 vdd a_n30123_n3051# 1.04fF
C970 a_n30483_7947# adsub_a2 1.43fF
C971 w_n28566_3528# a_n28791_3699# 0.72fF
C972 comp_b3 comp_b1 1.47fF
C973 w_n29898_n11250# a_n30330_n11313# 1.29fF
C974 gnd carry2 1.21fF
C975 w_n31473_n14760# and_oper_out1 0.19fF
C976 w_n26433_n9810# vdd 1.14fF
C977 w_n33912_n12969# D3 0.93fF
C978 gnd a_n29457_n10845# 0.80fF
C979 gnd comp_a1 5.67fF
C980 b2 a_n33822_n10638# 0.60fF
C981 a2 a0 0.82fF
C982 gnd a_n30330_n6516# 0.60fF
C983 w_n29178_135# vdd 1.86fF
C984 w_n29268_n2817# comp_a0 0.66fF
C985 vdd a_n30123_n10881# 1.04fF
C986 D0 b0 0.10fF
C987 vdd a_n35820_n11565# 0.60fF
C988 w_n28800_n4311# b3_not 0.93fF
C989 gnd and_a1 0.60fF
C990 D1 a_n28791_3699# 1.98fF
C991 w_n29547_n8685# vdd 2.02fF
C992 gnd adsub_b2 1.72fF
C993 w_n28566_5463# a_n28998_5400# 1.29fF
C994 vdd a_n33840_n1809# 0.60fF
C995 temp_more a_n28620_n5877# 0.80fF
C996 w_n29214_n5850# comp_b1 0.66fF
C997 w_n28566_3528# vdd 0.48fF
C998 a_n33840_n369# a3 0.60fF
C999 a_n30690_5400# adsub_b1 1.00fF
C1000 w_n30258_3528# a_n30483_3699# 0.72fF
C1001 w_n29448_3528# a_n30483_3897# 2.98fF
C1002 comp_b0 x2 0.41fF
C1003 comp_a2 x1 0.04fF
C1004 vdd comp_b0 2.34fF
C1005 w_n28737_n5787# temp_more 0.63fF
C1006 gnd a3 2.62fF
C1007 w_n29898_n4491# a_n30330_n4554# 1.29fF
C1008 w_n31941_n14400# a_n31851_n14373# 0.42fF
C1009 w_n33912_n9693# a_n33822_n9666# 0.42fF
C1010 w_n29268_n7146# vdd 1.62fF
C1011 a_n28998_9612# sum3 0.99fF
C1012 a_n29565_4599# a_n29637_4608# 1.62fF
C1013 w_n28404_n5085# a_n28323_n5166# 0.19fF
C1014 a2 a_n33840_n864# 0.60fF
C1015 w_n28566_5463# vdd 0.48fF
C1016 w_n33462_n3807# a_n33840_n3816# 2.17fF
C1017 adsub_b3 gnd 1.72fF
C1018 D1 vdd 2.17fF
C1019 a_n30483_10044# adsub_a3 1.43fF
C1020 a_n30330_n2187# comp_b1 2.31fF
C1021 adsub_a2 a_n29673_7947# 1.84fF
C1022 w_n28044_n5121# vdd 0.28fF
C1023 vdd a_n35820_n12033# 0.60fF
C1024 w_n33912_n14904# b2 0.93fF
C1025 w_n30258_5463# adsub_b1 1.86fF
C1026 comp_b1 comp_a0 0.40fF
C1027 w_n29178_135# a3_not 0.19fF
C1028 vdd a_n31851_n13896# 0.41fF
C1029 w_n28332_54# a_n28710_45# 2.17fF
C1030 AlessB_1 a_n27072_n891# 1.06fF
C1031 w_n28566_7578# vdd 0.48fF
C1032 a_n30483_3897# a_n29673_3699# 1.98fF
C1033 w_n33462_n2367# adsub_b3 0.19fF
C1034 comp_a0 a_n30123_n3249# 1.98fF
C1035 w_n29547_n3888# x3 0.23fF
C1036 w_n28260_n9846# a_n29457_n12141# 0.63fF
C1037 w_n26901_n9846# a_n26811_n9819# 0.42fF
C1038 w_n31941_n14796# vdd 0.28fF
C1039 w_n29547_n5850# x1 0.19fF
C1040 vdd w_n30258_9675# 0.48fF
C1041 comp_b0 a_n30330_n7812# 1.73fF
C1042 comp_b2 x2 0.90fF
C1043 w_n28332_n4275# vdd 1.14fF
C1044 w_n29898_n5436# comp_a2 1.86fF
C1045 vdd comp_b2 1.86fF
C1046 w_n29376_7236# a_n29286_7263# 0.42fF
C1047 gnd a2 2.48fF
C1048 comp_a1 a_n30123_n10881# 0.99fF
C1049 comp_a2 a_n30123_n5265# 1.98fF
C1050 w_n33930_n396# a_n33840_n369# 0.42fF
C1051 carry1 a_n29286_7263# 1.81fF
C1052 a0 D3 0.10fF
C1053 w_n29898_n7749# a_n30123_n7380# 1.20fF
C1054 a_n29637_8820# w_n29718_8919# 0.96fF
C1055 w_n29898_n10233# comp_b2 2.98fF
C1056 a_n30285_n7686# a_n30123_n7380# 0.99fF
C1057 b2 D2 0.12fF
C1058 comp_a2 a_n30123_n10062# 1.98fF
C1059 gnd adsub_a2 2.13fF
C1060 vdd b3 0.27fF
C1061 D b1 0.09fF
C1062 w_n31941_n13923# vdd 0.28fF
C1063 w_n29898_n10233# a_n30330_n10296# 1.29fF
C1064 x2 a_n28494_n1701# 0.06fF
C1065 gnd s1 2.01fF
C1066 a_n30690_7515# a_n30483_7947# 0.99fF
C1067 w_n29448_3528# a_n29673_3897# 1.20fF
C1068 adsub_a3 w_n29448_9675# 1.86fF
C1069 a_n29880_9612# a_n29673_10044# 0.99fF
C1070 w_n29898_n3420# vdd 0.48fF
C1071 w_n33444_n9657# comp_a0 0.19fF
C1072 x3 a_n28773_n7173# 1.16fF
C1073 w_n28566_7578# a_n28791_7749# 0.72fF
C1074 comp_b0 comp_a1 0.16fF
C1075 a_n29286_9360# w_n28908_9369# 2.17fF
C1076 D1 b1 0.58fF
C1077 b3 a_n33822_n10143# 0.60fF
C1078 comp_a3 x2 0.04fF
C1079 w_n27576_n5085# AmoreB_1 0.99fF
C1080 vdd comp_a3 2.20fF
C1081 gnd comp_b3 5.33fF
C1082 gnd and_b1 0.60fF
C1083 w_n35910_n12915# vdd 0.28fF
C1084 w_n33462_n3276# adsub_b1 0.19fF
C1085 comp_a0 a_n30123_n12177# 0.99fF
C1086 comp_b3 a_n30123_n8919# 1.27fF
C1087 adsub_a3 gnd 1.67fF
C1088 w_n29214_n1521# vdd 1.29fF
C1089 w_n29376_7236# a_n29673_7947# 0.93fF
C1090 a_n26811_n9819# equals_d 0.60fF
C1091 w_n29898_n162# a_n30330_n225# 1.29fF
C1092 w_n33912_n9162# D2 0.93fF
C1093 w_n33462_n1800# adsub_a0 0.19fF
C1094 a_n29673_7947# carry1 0.09fF
C1095 w_n29448_5463# a_n29880_5400# 1.29fF
C1096 w_n35442_n12465# vdd 1.86fF
C1097 comp_b3 a_n30330_n4554# 1.73fF
C1098 w_n33912_n12969# a_n33822_n12942# 0.42fF
C1099 D1 a_n30483_5634# 1.98fF
C1100 w_n29718_4707# a_n29637_4608# 0.96fF
C1101 w_n28044_n792# vdd 0.28fF
C1102 w_n33930_n2898# D 0.93fF
C1103 D a3 0.04fF
C1104 w_n28908_3222# a_n29565_2664# 0.19fF
C1105 w_n29718_2772# a_n29853_3078# 0.80fF
C1106 w_n27144_n792# AlessB 0.14fF
C1107 D1 adsub_b2 0.16fF
C1108 a0 b0 0.82fF
C1109 b3 b1 0.95fF
C1110 w_n33930_n1836# a_n33840_n1809# 0.42fF
C1111 w_n29898_n12546# comp_b0 2.98fF
C1112 w_n29547_n10647# vdd 2.02fF
C1113 comp_b2 comp_a1 0.70fF
C1114 comp_a2 comp_b1 0.85fF
C1115 gnd carry1 1.21fF
C1116 w_n29898_n1107# a_n30123_n738# 1.20fF
C1117 w_n28908_5157# a_n29286_5148# 2.17fF
C1118 x3 x2 0.27fF
C1119 vdd x3 4.30fF
C1120 D1 a3 0.07fF
C1121 w_n34488_n1134# vdd 2.54fF
C1122 w_n33930_n1836# D 0.93fF
C1123 a_n29880_5400# adsub_a1 1.05fF
C1124 w_n29898_n1107# comp_a2 3.54fF
C1125 w_n31941_n14796# and_a1 0.93fF
C1126 gnd D3 4.88fF
C1127 a_n30483_7947# a_n29880_7515# 1.60fF
C1128 s0_not s0 0.07fF
C1129 gnd a_n28998_9612# 0.60fF
C1130 w_n29547_n1521# a_n30123_n1755# 0.66fF
C1131 w_n29898_n2124# a_n30123_n1953# 0.72fF
C1132 w_n28260_n9846# vdd 11.96fF
C1133 gnd a_n30330_n2187# 0.60fF
C1134 D1 adsub_b3 0.16fF
C1135 w_n29547_441# vdd 2.02fF
C1136 gnd comp_a0 3.10fF
C1137 vdd adsub_b1 1.22fF
C1138 gnd a_n30483_5832# 0.74fF
C1139 w_n30402_3123# adsub_a0 0.93fF
C1140 comp_a3 comp_a1 1.18fF
C1141 a_n30330_n1170# a_n30123_n738# 0.99fF
C1142 vdd a_n33822_n10638# 0.60fF
C1143 D a2 0.04fF
C1144 w_n28800_n4311# a_n28710_n4284# 0.42fF
C1145 a_n30330_n1170# comp_a2 1.80fF
C1146 w_n33462_n3807# adsub_b0 0.19fF
C1147 w_n35442_n12024# D1 0.19fF
C1148 carry1 sum2 0.99fF
C1149 w_n29214_n1521# comp_a1 0.66fF
C1150 w_n29898_n9288# vdd 0.48fF
C1151 gnd a_n30690_7515# 0.60fF
C1152 a3 b3 0.82fF
C1153 w_n29898_n4491# comp_a3 1.86fF
C1154 w_n33930_n396# D 0.93fF
C1155 w_n29448_3528# vdd 0.48fF
C1156 w_n35442_n12024# a_n35820_n12033# 2.17fF
C1157 x3 a_n28224_n6030# 0.06fF
C1158 w_n30258_3528# a_n30483_3897# 1.20fF
C1159 adsub_b3 w_n30258_9675# 1.86fF
C1160 w_n28890_n7083# x3 0.84fF
C1161 vdd a_n33822_n8721# 0.60fF
C1162 D1 a2 0.07fF
C1163 gnd a_n29286_5148# 0.60fF
C1164 vdd a_n35820_n12888# 0.60fF
C1165 w_n33444_n9657# a_n33822_n9666# 2.17fF
C1166 w_n29547_n7146# vdd 1.95fF
C1167 vdd a_n30123_n7380# 1.04fF
C1168 vdd a_n30312_9297# 0.60fF
C1169 D1 adsub_a2 0.16fF
C1170 a0 a_n33822_n9666# 0.60fF
C1171 comp_b3 comp_b0 1.38fF
C1172 gnd AmoreB_0 1.07fF
C1173 w_n35910_n12060# s1_not 0.93fF
C1174 w_n29448_5463# vdd 0.48fF
C1175 and_a0 and_b3 0.54fF
C1176 gnd b0 3.09fF
C1177 a_n30483_10044# a_n29880_9612# 1.60fF
C1178 w_n29547_n10647# a_n29457_n10845# 0.19fF
C1179 w_n30402_7173# a_n30483_7947# 0.93fF
C1180 x2 a_n28773_n2844# 1.72fF
C1181 a_n29880_7515# a_n29673_7947# 0.99fF
C1182 w_n31473_n13887# and_oper_out3 0.19fF
C1183 vdd w_n29718_8919# 2.78fF
C1184 w_n28872_n5121# vdd 0.28fF
C1185 x3 comp_a1 0.04fF
C1186 w_n30258_5463# a_n30690_5400# 1.29fF
C1187 w_n29376_3186# D1 0.93fF
C1188 w_n29448_7578# vdd 0.48fF
C1189 a_n30483_3897# a_n29673_3897# 0.99fF
C1190 a_n33840_n1278# a1 0.60fF
C1191 D1 adsub_a3 0.09fF
C1192 a2 b3 0.82fF
C1193 comp_a0 a_n30123_n3051# 1.27fF
C1194 w_n26433_n9810# a_n26811_n9819# 2.17fF
C1195 w_n28260_n9846# a_n29457_n10845# 0.63fF
C1196 w_n33912_n14904# vdd 0.28fF
C1197 w_n29268_n2817# a0_not 0.19fF
C1198 a_n31851_n14373# and_b2 0.60fF
C1199 gnd a_n29673_5832# 1.02fF
C1200 vdd adsub_a1 1.81fF
C1201 w_n29178_n4194# vdd 1.86fF
C1202 gnd s0 1.81fF
C1203 comp_b2 a_n30123_n936# 1.98fF
C1204 w_n33930_n1305# a1 0.93fF
C1205 w_n28908_7272# a_n29565_6714# 0.19fF
C1206 w_n29718_6822# a_n29853_7128# 0.80fF
C1207 comp_a1 a_n30330_n11313# 0.60fF
C1208 w_n31941_n14796# and_b1 0.93fF
C1209 w_n33912_n11079# D2 0.93fF
C1210 gnd and_a0 0.95fF
C1211 w_n30258_7578# vdd 0.48fF
C1212 w_n33462_n360# a_n33840_n369# 2.17fF
C1213 comp_a2 a_n30123_n5067# 0.99fF
C1214 w_n29898_n7749# a_n30285_n7686# 1.86fF
C1215 vdd a_n29457_n8883# 1.60fF
C1216 a_n30330_n7812# a_n30123_n7380# 0.99fF
C1217 gnd a_n29880_7515# 0.60fF
C1218 comp_a2 a_n30123_n9864# 0.99fF
C1219 vdd a_n33840_n2376# 0.60fF
C1220 w_n31473_n13887# vdd 1.14fF
C1221 adsub_b1 a_n30483_5634# 1.98fF
C1222 comp_b3 comp_b2 1.59fF
C1223 w_n33912_n10170# b3 0.93fF
C1224 w_n33930_n3312# vdd 0.28fF
C1225 vdd D2 1.64fF
C1226 a_n29880_9612# w_n29448_9675# 1.29fF
C1227 a_n30483_10044# a_n29673_9846# 1.98fF
C1228 gnd comp_a2 6.23fF
C1229 w_n28737_n1458# comp_b1 0.63fF
C1230 a_n29853_9225# w_n29934_9306# 0.19fF
C1231 a_n30312_9297# w_n30402_9270# 0.42fF
C1232 w_n35910_n12915# s1 0.93fF
C1233 w_n35442_n12879# vdd 1.86fF
C1234 comp_b0 comp_a0 0.60fF
C1235 w_n29214_n5850# b1_not 0.19fF
C1236 w_n29547_n1521# vdd 1.95fF
C1237 w_n28404_n756# a_n28323_n837# 0.19fF
C1238 a_n28998_5400# carry0 2.85fF
C1239 w_n33930_n3843# D 0.93fF
C1240 comp_b3 a_n30330_n9351# 1.06fF
C1241 a_n29880_9612# gnd 0.60fF
C1242 w_n28566_7578# carry1 1.95fF
C1243 comp_a1 a_n30123_n1953# 1.98fF
C1244 a_n29673_7947# a_n28998_7515# 1.08fF
C1245 comp_a3 comp_b3 1.14fF
C1246 a_n33822_n15822# Gnd 6.54fF
C1247 and_oper_out0 Gnd 0.88fF
C1248 and_b0 Gnd 33.08fF
C1249 a_n31851_n15237# Gnd 6.54fF
C1250 a_n33822_n15291# Gnd 6.54fF
C1251 and_oper_out1 Gnd 0.88fF
C1252 and_b1 Gnd 31.42fF
C1253 a_n31851_n14769# Gnd 6.54fF
C1254 a_n33822_n14877# Gnd 6.54fF
C1255 and_oper_out2 Gnd 0.88fF
C1256 and_b2 Gnd 30.06fF
C1257 a_n31851_n14373# Gnd 6.54fF
C1258 a_n33822_n14382# Gnd 6.54fF
C1259 and_oper_out3 Gnd 0.88fF
C1260 and_b3 Gnd 30.52fF
C1261 a_n31851_n13896# Gnd 6.54fF
C1262 and_a0 Gnd 14.31fF
C1263 a_n33822_n13887# Gnd 6.54fF
C1264 and_a1 Gnd 12.22fF
C1265 a_n33822_n13356# Gnd 6.54fF
C1266 and_a2 Gnd 12.81fF
C1267 a_n33822_n12942# Gnd 6.54fF
C1268 a_n30123_n12375# Gnd 11.04fF
C1269 a_n30123_n12177# Gnd 16.56fF
C1270 a_n35820_n12888# Gnd 6.54fF
C1271 and_a3 Gnd 13.30fF
C1272 D3 Gnd 137.57fF
C1273 a_n33822_n12447# Gnd 6.54fF
C1274 a_n30330_n12609# Gnd 43.58fF
C1275 s1 Gnd 35.20fF
C1276 a_n35820_n12474# Gnd 6.54fF
C1277 a_n30123_n11079# Gnd 11.04fF
C1278 a_n30123_n10881# Gnd 16.56fF
C1279 a_n30330_n11313# Gnd 43.58fF
C1280 AequalsB Gnd 0.88fF
C1281 equals_d Gnd 1.86fF
C1282 k Gnd 16.19fF
C1283 a_n28152_n9828# Gnd 11.33fF
C1284 temp Gnd 2.34fF
C1285 a_n29457_n12141# Gnd 86.30fF
C1286 a_n29457_n10845# Gnd 58.33fF
C1287 a_n26811_n9819# Gnd 6.54fF
C1288 a_n29457_n9828# Gnd 48.53fF
C1289 a_n30123_n10062# Gnd 11.04fF
C1290 a_n30123_n9864# Gnd 16.56fF
C1291 a_n30330_n10296# Gnd 43.58fF
C1292 a_n29457_n8883# Gnd 64.10fF
C1293 a_n30123_n9117# Gnd 11.04fF
C1294 a_n30123_n8919# Gnd 16.56fF
C1295 a_n30330_n9351# Gnd 43.58fF
C1296 a_n29457_n7344# Gnd 0.88fF
C1297 a_n28773_n7173# Gnd 11.33fF
C1298 b0_not Gnd 7.18fF
C1299 a_n30123_n7578# Gnd 10.80fF
C1300 a_n30123_n7380# Gnd 16.56fF
C1301 a_n30285_n7686# Gnd 36.63fF
C1302 a_n30330_n7812# Gnd 43.58fF
C1303 a_n33822_n11583# Gnd 6.54fF
C1304 a_n33822_n11052# Gnd 6.54fF
C1305 a_n35820_n12033# Gnd 6.54fF
C1306 s0 Gnd 61.18fF
C1307 s1_not Gnd 11.65fF
C1308 s0_not Gnd 21.63fF
C1309 a_n35820_n11565# Gnd 6.54fF
C1310 a_n33822_n10638# Gnd 6.54fF
C1311 a_n33822_n10143# Gnd 6.54fF
C1312 a_n33822_n9666# Gnd 6.54fF
C1313 a_n33822_n9135# Gnd 6.54fF
C1314 a_n33822_n8721# Gnd 6.54fF
C1315 a_n28620_n5877# Gnd 11.33fF
C1316 temp_more Gnd 2.93fF
C1317 b1_not Gnd 8.22fF
C1318 a_n30123_n6282# Gnd 10.80fF
C1319 a_n30123_n6084# Gnd 16.56fF
C1320 a_n30330_n6516# Gnd 43.58fF
C1321 AmoreB Gnd 0.76fF
C1322 a_n27072_n5220# Gnd 5.08fF
C1323 AmoreB_0 Gnd 34.46fF
C1324 AmoreB_1 Gnd 20.13fF
C1325 AmoreB_2 Gnd 5.74fF
C1326 a_n27954_n5094# Gnd 6.40fF
C1327 a_n28323_n5166# Gnd 11.54fF
C1328 b2_not Gnd 9.42fF
C1329 a_n28782_n5094# Gnd 6.54fF
C1330 a_n30123_n5265# Gnd 10.80fF
C1331 a_n30123_n5067# Gnd 16.56fF
C1332 a_n30330_n5499# Gnd 43.58fF
C1333 AmoreB_3 Gnd 29.29fF
C1334 b3_not Gnd 10.81fF
C1335 a_n28710_n4284# Gnd 6.54fF
C1336 a_n30123_n4320# Gnd 10.80fF
C1337 a_n30123_n4122# Gnd 16.56fF
C1338 a_n30330_n4554# Gnd 43.58fF
C1339 x0 Gnd 0.88fF
C1340 a_n28773_n2844# Gnd 11.33fF
C1341 a0_not Gnd 7.18fF
C1342 a_n30123_n3249# Gnd 10.80fF
C1343 a_n30123_n3051# Gnd 16.56fF
C1344 comp_a0 Gnd 186.07fF
C1345 a_n30330_n3483# Gnd 43.58fF
C1346 x1 Gnd 36.32fF
C1347 a_n28620_n1548# Gnd 11.33fF
C1348 temp_less Gnd 2.93fF
C1349 a1_not Gnd 8.22fF
C1350 a_n30123_n1953# Gnd 10.80fF
C1351 a_n30123_n1755# Gnd 16.56fF
C1352 comp_b1 Gnd 416.68fF
C1353 comp_a1 Gnd 307.44fF
C1354 a_n30330_n2187# Gnd 43.58fF
C1355 AlessB Gnd 0.76fF
C1356 a_n27072_n891# Gnd 5.08fF
C1357 AlessB_0 Gnd 34.46fF
C1358 AlessB_1 Gnd 20.13fF
C1359 AlessB_2 Gnd 5.74fF
C1360 a_n27954_n765# Gnd 6.40fF
C1361 a_n28323_n837# Gnd 11.54fF
C1362 a2_not Gnd 9.42fF
C1363 a_n28782_n765# Gnd 6.54fF
C1364 x2 Gnd 51.94fF
C1365 a_n30123_n936# Gnd 10.80fF
C1366 a_n30123_n738# Gnd 16.56fF
C1367 D2 Gnd 152.21fF
C1368 a_n33822_n8226# Gnd 6.54fF
C1369 comp_b0 Gnd 337.58fF
C1370 b0 Gnd 87.79fF
C1371 a_n33840_n3816# Gnd 6.54fF
C1372 b1 Gnd 83.59fF
C1373 a_n33840_n3285# Gnd 6.54fF
C1374 b2 Gnd 75.06fF
C1375 a_n33840_n2871# Gnd 6.54fF
C1376 b3 Gnd 71.29fF
C1377 a_n33840_n2376# Gnd 6.54fF
C1378 a0 Gnd 91.84fF
C1379 a_n33840_n1809# Gnd 6.54fF
C1380 a1 Gnd 91.61fF
C1381 a_n33840_n1278# Gnd 6.54fF
C1382 a_n34407_n1233# Gnd 3.59fF
C1383 D0 Gnd 313.55fF
C1384 a_n33840_n864# Gnd 6.54fF
C1385 a2 Gnd 73.93fF
C1386 comp_b2 Gnd 327.30fF
C1387 comp_a2 Gnd 294.37fF
C1388 a_n30330_n1170# Gnd 43.58fF
C1389 a3 Gnd 71.74fF
C1390 D Gnd 106.69fF
C1391 AlessB_3 Gnd 29.29fF
C1392 a3_not Gnd 10.81fF
C1393 a_n28710_45# Gnd 6.54fF
C1394 x3 Gnd 73.38fF
C1395 a_n30123_9# Gnd 10.80fF
C1396 a_n30123_207# Gnd 16.56fF
C1397 a_n33840_n369# Gnd 6.54fF
C1398 comp_b3 Gnd 315.86fF
C1399 comp_a3 Gnd 375.69fF
C1400 a_n30330_n225# Gnd 43.58fF
C1401 a_n29637_2673# Gnd 3.38fF
C1402 a_n29565_2664# Gnd 26.35fF
C1403 a_n29286_3213# Gnd 6.13fF
C1404 a_n29853_3078# Gnd 13.17fF
C1405 a_n30312_3150# Gnd 6.26fF
C1406 a_n28791_3699# Gnd 10.80fF
C1407 sum0 Gnd 12.42fF
C1408 a_n28998_3465# Gnd 43.33fF
C1409 a_n29673_3699# Gnd 10.80fF
C1410 a_n29673_3897# Gnd 63.56fF
C1411 adsub_a0 Gnd 185.44fF
C1412 a_n29880_3465# Gnd 43.33fF
C1413 a_n30483_3699# Gnd 10.80fF
C1414 a_n30483_3897# Gnd 66.86fF
C1415 adsub_b0 Gnd 71.70fF
C1416 a_n30690_3465# Gnd 43.58fF
C1417 a_n29637_4608# Gnd 3.38fF
C1418 a_n29565_4599# Gnd 26.35fF
C1419 a_n29286_5148# Gnd 6.13fF
C1420 a_n29853_5013# Gnd 13.17fF
C1421 a_n30312_5085# Gnd 6.26fF
C1422 a_n28791_5634# Gnd 10.80fF
C1423 sum1 Gnd 12.42fF
C1424 carry0 Gnd 85.53fF
C1425 a_n28998_5400# Gnd 43.33fF
C1426 a_n29673_5634# Gnd 10.80fF
C1427 a_n29673_5832# Gnd 63.56fF
C1428 adsub_a1 Gnd 211.31fF
C1429 a_n29880_5400# Gnd 43.33fF
C1430 a_n30483_5634# Gnd 10.80fF
C1431 a_n30483_5832# Gnd 66.86fF
C1432 adsub_b1 Gnd 54.50fF
C1433 a_n30690_5400# Gnd 43.58fF
C1434 a_n29637_6723# Gnd 3.38fF
C1435 a_n29565_6714# Gnd 26.35fF
C1436 a_n29286_7263# Gnd 6.13fF
C1437 a_n29853_7128# Gnd 13.17fF
C1438 a_n30312_7200# Gnd 6.26fF
C1439 a_n28791_7749# Gnd 10.80fF
C1440 sum2 Gnd 12.42fF
C1441 carry1 Gnd 141.82fF
C1442 a_n28998_7515# Gnd 43.33fF
C1443 a_n29673_7749# Gnd 10.80fF
C1444 a_n29673_7947# Gnd 63.56fF
C1445 adsub_a2 Gnd 224.19fF
C1446 a_n29880_7515# Gnd 43.33fF
C1447 a_n30483_7749# Gnd 10.80fF
C1448 a_n30483_7947# Gnd 66.86fF
C1449 adsub_b2 Gnd 58.25fF
C1450 a_n30690_7515# Gnd 43.58fF
C1451 carry3 Gnd 0.76fF
C1452 a_n29637_8820# Gnd 3.38fF
C1453 a_n29565_8811# Gnd 26.35fF
C1454 a_n29286_9360# Gnd 6.13fF
C1455 a_n29853_9225# Gnd 13.17fF
C1456 a_n30312_9297# Gnd 6.26fF
C1457 a_n28791_9846# Gnd 10.80fF
C1458 sum3 Gnd 12.42fF
C1459 carry2 Gnd 131.59fF
C1460 a_n28998_9612# Gnd 43.33fF
C1461 a_n29673_9846# Gnd 10.80fF
C1462 a_n29673_10044# Gnd 63.56fF
C1463 vdd Gnd 1103.38fF
C1464 gnd Gnd 1551.22fF
C1465 adsub_a3 Gnd 245.84fF
C1466 a_n29880_9612# Gnd 43.33fF
C1467 a_n30483_9846# Gnd 10.80fF
C1468 a_n30483_10044# Gnd 66.86fF
C1469 adsub_b3 Gnd 61.87fF
C1470 D1 Gnd 980.84fF
C1471 a_n30690_9612# Gnd 43.58fF
C1472 w_n33912_n15849# Gnd 29.29fF
C1473 w_n33444_n15813# Gnd 28.07fF
C1474 w_n31941_n15264# Gnd 29.29fF
C1475 w_n33912_n15318# Gnd 29.29fF
C1476 w_n33444_n15282# Gnd 28.07fF
C1477 w_n31473_n15228# Gnd 28.07fF
C1478 w_n31941_n14796# Gnd 29.29fF
C1479 w_n33912_n14904# Gnd 29.29fF
C1480 w_n33444_n14868# Gnd 28.07fF
C1481 w_n31473_n14760# Gnd 28.07fF
C1482 w_n31941_n14400# Gnd 29.29fF
C1483 w_n33912_n14409# Gnd 29.29fF
C1484 w_n31473_n14364# Gnd 28.07fF
C1485 w_n33444_n14373# Gnd 28.07fF
C1486 w_n31941_n13923# Gnd 29.29fF
C1487 w_n31473_n13887# Gnd 28.07fF
C1488 w_n33912_n13914# Gnd 29.29fF
C1489 w_n33444_n13878# Gnd 28.07fF
C1490 w_n33912_n13383# Gnd 29.29fF
C1491 w_n33444_n13347# Gnd 28.07fF
C1492 w_n33912_n12969# Gnd 29.29fF
C1493 w_n33444_n12933# Gnd 28.07fF
C1494 w_n35910_n12915# Gnd 29.29fF
C1495 w_n35442_n12879# Gnd 28.07fF
C1496 w_n29547_n11943# Gnd 26.52fF
C1497 w_n29898_n12546# Gnd 73.22fF
C1498 w_n33912_n12474# Gnd 29.29fF
C1499 w_n35910_n12501# Gnd 29.29fF
C1500 w_n36234_n12420# Gnd 28.47fF
C1501 w_n33444_n12438# Gnd 28.07fF
C1502 w_n35442_n12465# Gnd 28.07fF
C1503 w_n35910_n12060# Gnd 29.29fF
C1504 w_n36243_n12096# Gnd 24.41fF
C1505 w_n35442_n12024# Gnd 28.07fF
C1506 w_n33912_n11610# Gnd 29.29fF
C1507 w_n33444_n11574# Gnd 28.07fF
C1508 w_n35910_n11592# Gnd 29.29fF
C1509 w_n35442_n11556# Gnd 28.07fF
C1510 w_n29547_n10647# Gnd 26.36fF
C1511 w_n29898_n11250# Gnd 73.22fF
C1512 w_n33912_n11079# Gnd 29.29fF
C1513 w_n33444_n11043# Gnd 28.07fF
C1514 w_n33912_n10665# Gnd 29.29fF
C1515 w_n33444_n10629# Gnd 28.07fF
C1516 w_n26901_n9846# Gnd 29.29fF
C1517 w_n26433_n9810# Gnd 28.07fF
C1518 w_n28260_n9846# Gnd 161.09fF
C1519 w_n29547_n9630# Gnd 26.36fF
C1520 w_n29898_n10233# Gnd 73.22fF
C1521 w_n33912_n10170# Gnd 29.29fF
C1522 w_n33444_n10134# Gnd 28.07fF
C1523 w_n33912_n9693# Gnd 29.29fF
C1524 w_n33444_n9657# Gnd 28.07fF
C1525 w_n29547_n8685# Gnd 26.36fF
C1526 w_n29898_n9288# Gnd 73.22fF
C1527 w_n33912_n9162# Gnd 29.29fF
C1528 w_n33444_n9126# Gnd 28.07fF
C1529 w_n33912_n8748# Gnd 29.29fF
C1530 w_n33444_n8712# Gnd 28.07fF
C1531 w_n33912_n8253# Gnd 29.29fF
C1532 w_n33444_n8217# Gnd 28.07fF
C1533 w_n29268_n7146# Gnd 26.36fF
C1534 w_n29547_n7146# Gnd 25.95fF
C1535 w_n29898_n7749# Gnd 73.22fF
C1536 w_n28890_n7083# Gnd 161.33fF
C1537 w_n29214_n5850# Gnd 26.36fF
C1538 w_n29547_n5850# Gnd 25.95fF
C1539 w_n29898_n6453# Gnd 73.22fF
C1540 w_n28737_n5787# Gnd 161.33fF
C1541 w_n28044_n5121# Gnd 29.29fF
C1542 w_n28872_n5121# Gnd 29.29fF
C1543 w_n27576_n5085# Gnd 95.92fF
C1544 w_n28404_n5085# Gnd 28.07fF
C1545 w_n29205_n5004# Gnd 26.52fF
C1546 w_n29547_n4833# Gnd 26.36fF
C1547 w_n29898_n5436# Gnd 73.22fF
C1548 w_n28800_n4311# Gnd 29.29fF
C1549 w_n28332_n4275# Gnd 28.07fF
C1550 w_n29178_n4194# Gnd 26.36fF
C1551 w_n29547_n3888# Gnd 26.36fF
C1552 w_n29898_n4491# Gnd 73.22fF
C1553 w_n33930_n3843# Gnd 29.29fF
C1554 w_n33462_n3807# Gnd 28.07fF
C1555 w_n29268_n2817# Gnd 26.36fF
C1556 w_n29547_n2817# Gnd 25.95fF
C1557 w_n29898_n3420# Gnd 73.22fF
C1558 w_n33930_n3312# Gnd 29.29fF
C1559 w_n33462_n3276# Gnd 28.07fF
C1560 w_n33930_n2898# Gnd 29.29fF
C1561 w_n28890_n2754# Gnd 161.33fF
C1562 w_n33462_n2862# Gnd 28.07fF
C1563 w_n33930_n2403# Gnd 29.29fF
C1564 w_n33462_n2367# Gnd 28.07fF
C1565 w_n29214_n1521# Gnd 26.36fF
C1566 w_n29547_n1521# Gnd 25.95fF
C1567 w_n29898_n2124# Gnd 73.22fF
C1568 w_n33930_n1836# Gnd 29.29fF
C1569 w_n33462_n1800# Gnd 28.07fF
C1570 w_n28737_n1458# Gnd 161.33fF
C1571 w_n33930_n1305# Gnd 29.29fF
C1572 w_n27144_n792# Gnd 62.16fF
C1573 w_n28044_n792# Gnd 29.29fF
C1574 w_n28872_n792# Gnd 29.29fF
C1575 w_n27576_n756# Gnd 28.07fF
C1576 w_n28404_n756# Gnd 28.07fF
C1577 w_n29205_n675# Gnd 26.52fF
C1578 w_n29547_n504# Gnd 26.36fF
C1579 w_n29898_n1107# Gnd 73.22fF
C1580 w_n33462_n1269# Gnd 28.07fF
C1581 w_n34488_n1134# Gnd 41.25fF
C1582 w_n33930_n891# Gnd 29.29fF
C1583 w_n33462_n855# Gnd 28.07fF
C1584 w_n33930_n396# Gnd 29.29fF
C1585 w_n33462_n360# Gnd 28.07fF
C1586 w_n28800_18# Gnd 29.29fF
C1587 w_n28332_54# Gnd 28.07fF
C1588 w_n29178_135# Gnd 26.36fF
C1589 w_n29547_441# Gnd 26.36fF
C1590 w_n29898_n162# Gnd 73.22fF
C1591 w_n29718_2772# Gnd 41.25fF
C1592 w_n29376_3186# Gnd 29.29fF
C1593 w_n30402_3123# Gnd 29.29fF
C1594 w_n29934_3159# Gnd 28.07fF
C1595 w_n28908_3222# Gnd 28.07fF
C1596 w_n28566_3528# Gnd 73.22fF
C1597 w_n29448_3528# Gnd 73.22fF
C1598 w_n30258_3528# Gnd 73.22fF
C1599 w_n29718_4707# Gnd 41.25fF
C1600 w_n29376_5121# Gnd 29.29fF
C1601 w_n30402_5058# Gnd 29.29fF
C1602 w_n29934_5094# Gnd 28.07fF
C1603 w_n28908_5157# Gnd 28.07fF
C1604 w_n28566_5463# Gnd 73.22fF
C1605 w_n29448_5463# Gnd 73.22fF
C1606 w_n30258_5463# Gnd 73.22fF
C1607 w_n29718_6822# Gnd 41.25fF
C1608 w_n29376_7236# Gnd 29.29fF
C1609 w_n30402_7173# Gnd 29.29fF
C1610 w_n29934_7209# Gnd 28.07fF
C1611 w_n28908_7272# Gnd 28.07fF
C1612 w_n28566_7578# Gnd 73.22fF
C1613 w_n29448_7578# Gnd 73.22fF
C1614 w_n30258_7578# Gnd 73.22fF
C1615 w_n29718_8919# Gnd 41.25fF
C1616 w_n29376_9333# Gnd 29.29fF
C1617 w_n30402_9270# Gnd 29.29fF
C1618 w_n29934_9306# Gnd 28.07fF
C1619 w_n28908_9369# Gnd 28.07fF
C1620 w_n28566_9675# Gnd 73.22fF
C1621 w_n29448_9675# Gnd 73.22fF
C1622 w_n30258_9675# Gnd 73.22fF
